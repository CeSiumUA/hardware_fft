��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�[�ק���dI ��Y�l�BY�nyWE��:�0`��}�a��R����1.�_E}�>���ۺ�FI7 D��5�1k�.�@GdQ���(3J��U���6��ɒa���6?Q0�^B���DD��H�����u�Q-�l��ݵC�=������s�k���&p���e<��x�h�-��4���;�f��W�6���w.�[�0�*�ďQD��"D�?Gd/�/�[M�@�k��h,�e}�|�/�6�4%5E����-�G�nec%;Ԧ_?fTZs*�K﷑n $���kN0�?�ψ?����茇h���V���=o�Q(͝3�U�dd�f���;V��/���.�_|��ܡmm��p4x*+��K��o߭(l�JhtP��C�i��m���n�gR�	S�n�����ȏQSq�~	��d�e��Q����O�+�'c�{W���l�`-9�o/��\椋��tBxW�h�F���{�#�Zh�������Y)o�O��� u4ب���
aL�u}��晣;t���2Jl{�Cj{�h���A���J��7��p�{e�:�(m%V9��+��hVu�S<A� >|�{�y+%W}.�n�t(�.�3�$p2�3�ᛸ��ݫ�ǐJB�2���	(T^ ��8\l�p`��7R���V0u��7,&}0�ܤ$�U	&�`�1�W���(���N�|����2H<��7�P��
K�Ef�o�/Z����Z��w��\�ǫ�]��W���#20�lߙ�I����ta�I��(o���&Ե�t�k%�.�[�0����h�	��rW��h7��=88~Z4� �~�vۆ�mP��~]�Q�� ��f��;e��CRlv1|ӷ���P!���É��}�Dr7�a���^4�@V1q�#�*�Ed~�׈�ی-��|青}���j�yH��'ZÉ+e�[C��=s���)�g>>�VG��W���\���稌8�܍1��P���v9K��N�
T:��-�_���V�������L���d#�GDo���C�a3�K�����x���^1��tD�������<�����c��J�5<�R�L���`���M�w߈Hqś�;�[
��rŵ'|�b/rY��$��	��2�Y�MC�L$>Ғ�vE�N;�J2�����8�	��X���\!0}z4=���Pe�M %ƞ�	�U�T����[ᭋ�@��֢ G~x ��������諢��,��=�<%�˄����^sW2\R�;$ �,ub���M�
���?; ������0��^�g�&��k�#�>�?1�Yb��*���fs�2���߯�i:ǯ�'�'d���]*��~<�}��A�%N��{A��:@�*����~l��S6#޼_������=�N��x��Z��n�+T�����V�k�%h��nY�tA�"�*�ȈU##���ز`������D�Hv����L7����s7���3 �̸���LҾ��E.��FL:�J�A�43��3����J�w)ՃA7�'#)�3�'K+�x����s*đob̗Y���7ԯ��`�xB��)��v�7wu�5��u<�-�J�
�T�aIa�����`�m�?���������8��%6��λI��� "����h�(������.~�)A�t�k=��y��d��4\¬�
�3u��!v��W����~���)�ioĨB�uL{�шE�xFW�Ѫz�n�'{�b"y//�R	�/{a}B,��;�(v�@ʿت�WB]��?;����3���s�=�켅�H(
Q����b�����1�:�W�P�Ys\l����=b��<�7�f�/Q���S��>���O3�oTZ�_�Y��L�k@u͌�$4��);F����)��@�s/:�x�����M����ʡ�jp&�8Rb��_���y@w�9�X��P<S+�R.Ŷ�m���3�{�A�����%�aΡ���0�bUƹ���"�Ǧ{h$�/#�a{U-2)+[��r�,��{Ľ�9/3�{g�m����$��Z�o�.���6�ň.��A�}`��l��^nkT1Bv����*���f�Z��m������8S <���?"��Q`T�u�|�{�����9�:*��ک����T觝�Z.1�$)�^p��!�q��/��(��5*gŨ�K��H�4��A}H�����6����4U���@���5e��u��w-�q	�t�/x����&q��LG퉐1���X|�1P�'Ѐ{�l����<i0����`�&���E#7�aj����O�=_k>�̌p�vCz{�L@��M����+��A��p�(#!%p�y�Ƶ��[�s"@V�=��q��f�ƞ����{���ӽ�%���!���Sc����Ҏ��ڬQ��/u�f��) `�Zs��'f��{��j�q��='�~ `�p�6�����W����	(9D�30(D����I�����b޶x:�O�p{ҥJhO_�w�y݀�W{�0�(D��nr5P�w��	G�2[a�QY�or�Q$�+�g�,�S�	�/i勒�~<kH��Fy��t}�,b����H'T?WqW#>cvX�ܤX�{[٧Z뉰T]�kv� U��pˈ�^B��' @��Ŋ�C��?2�t/����ڃ�v�
Q��m��(���Y��R@3,��$�3e$�%P*�Y�˳O'��>4,;�ZHUyUMhs��T������?��u��h���)c�a�����H�Q�M���Af��*+ĭt[Suj��f��b ]T����L���T�k̾�][BT�m��1�E7��=EӀ껹a�!��(��@���"Ej�Y�0��_/��'��ͬ�"�7j�9��}��mGp�:}�Q��`G?n��7����Ϻ9W��\���3�������-�Q
D�HȊ���4�����xw/�٠KV|�G�&u���;�w���nL�v�S���a�ѡX�6��8|���ǇԳ��'������(�U��N��p�-���<���o&�w�����K� ��F3tԺ-Zy��2�sه���Q+��	�=]��Pp'���AV��ϥ��N�^(��㥫�
	�濧d����)��<�v �(C*���mT�^=� �����U�y$1���j6���ϾQ���DD�u�F�1n1ߚnWp��pO�� �5�`�7��g�e�ږ�oQ�u�p]����PW�uT	)>�Ĵl�� �/!�7�5F�Єz�F7�o���$r��P��U`-�{�Db H�Ϻ����c�b���P�M��"~>����;0���NA������:}�PI.�xQ�v2^���o�-��sh���y��FKis�����<�L�^���� ��X�Ƙh'�9\�R�b.��qg,|�en�����+5<d�Q�H����5���Xl�K�����:N�u8񙰳���CB�cʅ����}�\��#qr�8M�֎�����FLgkt $��s�.fB㭇�/�g�%��2H�W�"f��aɣ{eg'z�D��'��yK��#���_Y/�2c��$