��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B�� L���,F��+*2 ���n��E�L�n��R���DG���:L��$۶7�V[)3�����כCmO�"��Wߊp���(��DU�����`��N�s$������EK��N)��s�����q�"�l�bJ�ٕ"=wH�_t� �гW~�9�!�1�5�E�߯9����4+K0�厕1�� �m���=fҵ�*��g|��,˧<���Y������R�T\a�T����WV��� )�xӛϒo���혛�P��g����;dF�SGܶA�%;�3�2�]�-�+N��s(}^5�4����������^��ꗑS�#6.��Y�k�h-�|�v�~�Li[�xg��KIXX� $����7q�h�0*�Ah���L+��^K#��װ�M�yJI|)l-ř��w��py��@�^��0�}�)�Įچ�ps�#���*�`��_�Cl��C�h]���u@�H!JE� �~N��>�9Q�=�K����g�	ر�-c�`'��B��>�q���!r�J�h�p�L6�LA{�f?O�e�G��n��ȹ �Y�^�nAG2�N��R�W�u�$������G��8ǰb�M|M��^dG��)������1Z02��T�v?���̨pE���tD6��ye>`UPP���-�����뿆u�W+��x�Z�[�>,��������E�j�j	�9sʣ�S��6Pm�@��}_�YZ���J:����ͶD�GBVW��87�+��g��a�$��W�l�����Uj��6zD��e���A�H�Ʀ���^��=Fp�}�@����� ��?,y�P�Z���yO�8kx�\�l(?'��`N��������O&<v��[W�/S*H��]�#n�����4G���m�Gd�h��5����i�_Q�Q�#�\˞��Hv�o�^D�F["�vE� �É=�(��8g豈?RK(�8���E�=���䳕��ASW��ڿ�f!�-Y� g]�'NmB���w�Q�,���͕k�U4��@�q�e��O���D5���ܑX�[!z):����+�(1 ��]Y����}����D�kmp)�:�I��!���;s �t���~BQ�=!l`v�|흨��y��:����
��P�)P)���X�b���潢��}C/�
��L��t�����{2�;��R%
!$X`i�ƿj����Q)��/3���X��{�y�@򰸙v��g���O���<F��^�����ni5�y,$p�����L/��̦д6~����Y'��_�������rX���b��
n�{n�j�l�� �ϥ>���s�t�Pwת©R�5�מ\�d@�������(�C�K�o���W����([��ٞ�D`%���_� ��Q�(Bnͬ���B&�_=�F6�c�Vl�q�=��������6�rUO^��Y��4\��}�~\�m�w{V��'����߬��^���jco��/�Zv�|c�yCf�2J	�7�i$����2��>���Q��L�N �uSg�,�CB�\W�x���;8#�:���ި��	a@��䃥�p_$�> tzቓ�z�.=L��A��G�d%�n�;��j�������:�6��4��\\^{¡�bɓ�*��w��ߓ5��ب����v�ލ��Qh_#;쳕J�ޱB�cM)��M-��p��b��C�!��T6&S$c,s�����J$(Z�.]�[����� �<����bN�<S=	-��#�<�n����jh	����OJ��Nq�'�S�Uq�qmצ�Rǟ�L��;�^9��68�^͛ޫd�^��'��<k9�tw�\�*��~i�~T�!�SΦ��;�]�_[>O�6Ni�4��,5�?4<R�O�f�Ã�W�������H]���L�s�.���	P�z�|D�!��8/�D��MtH�y�Xm�_����7fu�,�v�g��J[���}7?f1�X�j��k�=�c�c�d� ����2��f!N� ^�+��?��2`��Ʒ2�S[���bӿ��1|[Y�ծ�Bf%ˀ�c��O8��P3�!2���B]ڕ�j���� h�23�>���3����*Ȟ��� ������1��X+o.gPO)�vm4��w#P�@�t�p��H�=����n�?�p�m�>C��@�/����_�=�#��|�jm��Ü�4�2%Ѭ��ݸ�