��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w���>��!S��'ho)�mRv��� �=ß��;��!�����=-�F�'��-��$N�9_Ta}u�~-����jL�(�s{1�Cy������[9o{':�����C� \�(��Z�`U����;į�n	��o:�5Y��uU�b�Q�Ć�����@Ml>mo؂�R4V�ڨ��퓌�r!���ԇ��T*��N�f-���剪���2�)�����}�htܤ3ǔ_�ΖzV~ݰ���OB_g+B��$���퐖��ʷ��Mh\4�w�ҵ��8�ęQ�,��\�Y^�!@�ǄX�l�����l��%?a������Z	��vUN�J���ý�0-�j��8�8�}�X��O��]&�烾U)�k�,���~�״}_��pEV�4�����`���5.�M��%e �:�L� ?c��h��/��k�qfvF8VSI�f�6z���Z%�A�SLu.�����f�0لUP���K�5����H�dzc���6 ��uҙ<-���3�B߾ �	���0�p=�ݰ/r���l^�IkH�g3gn?���>���&v�2�\B��Cã�K&wS��;&���?�Wp5I+H,��������s�㈕��k��d�� N�������a��� �M��ygǆ���s��50u�/��ҩ��]����oV������g�0j���ҝ���hԉ�����j���ѧ��9�\cyes���h��nIv�j&�J��W:'Ǹ��/�\!�`9��%��E�QR9O���.�S���$u�����4/����Ct���
R��K&��~ɔ�2B=0��NRw:[�>�xq�+���"^I���)3��%��ۏ���T�r�t1�k'�N��ż���9"�b#H� �&T��Hc%,=n�G�s��V��b��47���!��B?�(g�==��d%ynp@�u���Oud��G��K�Rg[g�*�T��2��*�ۥ:�މ���`�1�-=���)���C��q�5?"/��5�zi��R��:,�uN��:.r.�fYE�^���I��d����m�HW=�&n��Z�^�}�q5NΡ �^�f��(�u�4��2�,�0��C�)�@ ���N��w
�6���|>Zm�4�g,���Wڳz��o��H��P�6B��K�����FɎkӔn�jf%�P@��|�6i�7 �RE����Z����[�]b����טs%m�v�w�����!(,�ٓVG�@���n�(N�d)ia��Mr���WZ!���|�#�Ԑ�����%��:�\��\�������I�s��\C��İ��Ƿ��:�'����`ByiqXͤ|l��m�Eǋ}�&$�ֽ誻�x,+�w�*z�w�$g���B7 �)Ti���S�������϶C*ő�/fV2�n+?=KP߀]�x�w�CJ�����$�1�-m4U[�l�Y�,fs���5g9�f V���7��)������BM��D�Qv�X����3u �q����f9�Qd�<Cx��{�\�����>[�X�?��9fL �2���I;_�H`�hNZ{����JlQ��u�宭Wף�91U/_A�!���oփ;����h�I�S��DO"�>�c�ሼօ���m-E�,��U�9!���&Ŋ�c:Qd�?X�1�>�a�ʟ�Sξ�pjA̳�@1��@Vg����04:Q^8Ά��z6����5�S�,r���bM쯣�$3�5����m��Eb�l~�@�f #U�P���ݎ ���q�6���� g�Xs넏�<�+�+���4!���ɽޝ� D��ܞ���`<8~�ϛ3��X����0u��}v���n�Rxm�]��Ğ�C~�X�~�R�����{�oi`�˭r��.��edӗ���w�b_Xz�b)�&�DN����B�'@;��E	̬�+ڪ�:	�����Y��i��1�<D��Zo��-����ެ	F\�Ǘ\-��M��jl�?Z~LR	�f����e��W1aU��s9�m^�9�ܞ2e��䎝�%��l,AHd��L��jv.ų�2�P����B�������D�hJ�Yt������q�nkѸͭ�m�ஷ�h���_�Lb���>ҽ#�2�����6���J�bF� �H� �r�H����gey�5}�\�/�q�ĭ�JB�A���_���Ы�7�qa% �V[BY��v��VIE��w���E����t�`5ū��[���N�#K1����\�hk�5r�'�H������?5]���K"�~��.�5��@����g���4gdx�);��������7'�G��9���K('��:�t'�f��Y��r'�=�����A+o����j���4�_��_咨`e�j�楏��$Lr�e�����I��7���B���#}���v�9{��W-�z[:O��V�PW�gQz��&NĪ���ǁ\�;�EK�LB������p���d�i�	�񈮎a��D[��o�@8�i�`�L��o����j�v|9+m�x�P��KT9���ӬF�������?^�°q̉o��!7"�/�l��+~�1�3�F�㠢���'�Ͻ�t� ���PNriE���]�V;�y�ްPK<��'K� ̣�~$�L�C�u��Y�NWp-J}�i O
1
�*�����M�"�E�6�XgPH�Y�8�#n��Ģ��<S��KbY�(�(��~�"� �g��l����+z�	�Be�DN6�:wr�A[��0|�x|0�t��[p4dS����RL���:?�׌5����nU��Y~]��8����߸���[��B��5q�w�\}����b����~�RD&
��p�R(�1�#{�����nfR����e֤��o�l����B�]@�q�޸
�x�t���#[ݸoy�����C�CW�jb$������UrT�y]h���0�P�&�s��g8ӽV�n#���oX10J\�q �W����.�|Y���J�O��*���p�-�����M��xe5p�wy=���=�������E���ɋI32���\����xê��"K<��3��L�۸��Fz?% �T�ӏn hXmN���;��Ip�%O6���D��@D��~��qv�́�4�O� 3w#���B��P�5�0���ީ��>�W�m(��2K�e��y���1 ��|�%�u�������p��V���Cb��}�Y�װנ\��yNh��ݨ�s<,iN�rx矞�}�!�JqO��B� Ծ��b��3��J:�V�X��y��g���Pou��y���YLur[`�����&\�0�f�T�#���tpÓ���ψ�h�����#ﾎ�&�f�U9Jp�t�)~�l�0�"�ϧ�=@�07� E���f��
ơ�L�����L��'Ҋ�i�W~!�#�9�E����d��:�k�L֨7�=�����z�5"��}�BA�x��$�kP5M���KE�)��(�pK�۔��%Nc���ٺ�
��odѝf艌��n���� 'Ks���T�:>�G�D���2tT!�T^�s�ɝ63k��wN�����Ԣ`Q̘>n}SJ��h�6"�R�������`�2�X�L��/��xK�>�):X
���0��.���Fϴʻ����4)�l7k���__n�||��Jo��?�m<�\�W����>y�V&l ]e%*/"�W�
`���ԢC��h� ���^�AT�	Vvpܬ;�F��).�ՙSVw e��w��y")�Ԙy��3�I�F7y8&��^������������ڵ��̰�(\/����3�v3�l��bLT�:��)�,��=ן~��n�e�{a;;N(fB_)|�ގC��8�����T� ���k+�q�kc�DY̢&���5G��<Ϛ"�~����C�bW?��f<���SA��qV�+U�yR�`�������&Cx����kGa��zK�xNƁR�@Ճ]4�wv�j*�6֖�g>+=*���jc�����`�W�B�mWJ�[j��l�<�CJ��Ū#������f�U�Zm�a�8�wC,<x)���+U@!#�l	�M�I,-���vw����/L<"pw���Ҥ8�@fYڃ,���~�O77�����f�̸Z0���d��]�̯��R���eKo~�L�B����:�S��믂!4'���N��X�w�H�t�+>�-��Y+Q�N�%IP!��rQOEF���&ؾ"�e�������G�:�Ν)8~���fe���Ӑ�+���n���Q��Ϧ�DY�����)\���0���M�в�xA n���#�� ��Qd_�!���oT�8�f����7�y�)�{�^_�������رLy�c6���w�Zw$ �(�jYxg"4���[��~ɾQ��&M��$��ނ��Z���5P�Yp���! �H �]���P��TQ��1�����D���@�)�l%U��;�sV�)^�%LV ��3�{����B���t�ڒR�Us8���ǭ���� �;Ja+s�a�8z�~�%m�8���Z8�g��5�aaս��N_Xb:�l�t��'�=��dI	�)`JA�y*��!�e�#Ć��KO�&m���.b���tR�?ߛ*hp��@��)^�"���j,�''����p�Q����ƥگ*��ü�_Y(I�g���-lԦ`�M�j	��h+�t���x�����/-����B~օ�ٸvߩ��+�h�sA6��d��F����AhU���_kh�J%�][�'���}��g����r�UI��l�5bgQS3�$��2�jܥ�S���%��/�w�`J ��8<�Ɓp�3·{�X����,�K��18�Q�8�Gj�U"�x��� 7g�f/��ޛ*�әy�`�Aw+���JS'��(,m���6i���@�����F�n���g�*�㋇ V�<pnb�����nL�}��zǥ�"P=N���YW�b���$ݙ�~=K�T�����+��zv[9F��/R����*�����O�	�� +ܻ�����P�?!����&��8c���6�)6�_�6�L��!e�x$��:2;�6�E��M{���0P�I�,_�/{�����q(s��修�=���Be+���Xs�z��T��yFҾ% ��+[�^���a%f�b��8�}�"u!=~��>�;�(A��v>:�ߑ5��\e&�D2
t�S/y���^��/xY[��r\7��ɴ<%��	��o� J@�u]N�zg:���c����AU���,�i$����^���~�Ci��_:����gvw3��4l�"��p¹����<@s�/��h�$�y��M�*|��@��ݮԈ|ܐB2~�J�"�C���0���/���V��2Qئ�FmV*9�X�1�;���d�}�;K���E
���[��h���20�*�ǒ�Y*�b#���+08?�̣��������-�9�\�G�̈��ŷ!�-Fwy��AMȩ�`KO�qŚZ�P�7s4���p?8Y��zat@ۂ���@ք�\�Vw�����H� yϧ�R��FMV�c�B0��E<o.���xV����DOVF]�Ӡ���?!zAq�Zp�c�����jkX�3	��`���d	���Uh�N`)[#�䷹�5h����^��0<��ں��'8����F�>B�����$%�v2�j+���fʹ��v�75_�k�2�:-����Y;���"����P_tٯ��BL �ѕ	��BY�s�m$ ÆE�z�&\0ÝHk�������R,��܄HD1^g]�m����'u���UE��"�D�x� &m]^/�O3��z�f��`V���47�|&;n��d�5Ķ� ���+S����@_O��Ao ,��3 3z�]�:Fc�nf�*	i\���Om
cK�@t��]�I:\�(���X��vb�����1�W�L��CP:�\>��3��떵y�e�ip�r���E�OU�)!�؃2�򞫻:�҈B�O�m:j&�P�9N&K 0�Yf^2�p<.8P����$�����#U�k�:n'h���<�Mn�̓�įo5̡8<�sO�?�*��o8��WC9P�Р$��ͫ�y+��v	X	���4�5�n�f�Z��d��;Nӿ� 1��D┪)���