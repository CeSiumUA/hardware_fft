��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c��P��OK��F��/�v�<j�}.[�6�Ć��6 �������t'���5��(n&�4��ҪX��Zr����r36k%ѾW0U&��:t�)�s��C-Uz�#T84�^$:t�(�}�N ����&SYI�X�" ����Y��B(R����������'A1���n��8C[����j�����·7��U���L����k��ܻL>b�����ʊ�)R��DJ:
*ř�ŉ��P�g_���1���d�	ȥ� ���>-�u���lu��Uš[��-x�Qeۜg��[ц��
͝S�-Q\+?��l�3���*5sf �.P��:}l��񿙁󨀭����`�����5��2�� X�
ڄ%&���U���خQ�$�T���e�۹�
��ѭ��,���?[����+7Lb)�0�f��o���@��:�c�����ͯ
�tR*s��{�ah�0�p���ͣ|��f��M		��7G!�C��Hd����ױ�:��H@�����-���r:	6B�E�������C�� BR�Z9Kh.6�\�wH�8|A�P��}�wFH�sc/1�zm:���c|�0��,����S������Z�LB�k������0�b��0Mu�g��'������K^�^tk�Z���)6�
���Z�k(7���&5E����l�����ь[I�9w���TH>w1��?=7\P $�K\��_�{1~��0������(�ּ� ڼ��@�b�0a��?���=�y#gc{�E������mDt�sF�*�WJ-�"wuw���E�+�%�����|��ɗ����&@$�9���@Y!Xgy�Ս@���}J��Q��ٻ��ku�O���g�gN �u��)nC��^\;R�Q#)��i�6M�b�a�[���*4f�ׇ�JT�XD���e�L�Ki{����q�5����3+�Q��;�Ѭ��|�����L���#I�!H.[b�c�G��ƺ%oj5�����i��o܊r�o�C�$�y��,�D:�W��Q8���H�pqX�ॲ�y����r,)�34?�TǧA�̅��t�Ȯ`Ϩ�t�g&�� ���']�2O�.�|o�ϼ`vo�+N�F�I��?v*�o/f#ȩ+��@���U� wu�A�'v~��V1�Q�\՚����ȡ�-h�=e��`½��u�L9���9��b+�拎c�J�#Sa�dX�0#h`�ct�M�P0�r!Xed�F�<�z���ޫ��?��7�y��x�@2��u��$HڻE����y���	�hSz��ҫ�>�O)ߊdlR���v����������T�$�����8t	��΃���h���~{t���m`�+��~H��=�&�q)�-͡V��͵���b��.+�ė�J��Qw-yJ��9}�F�ۣ�\�^��$�-��	�.p�P�����m��E�v��"xV��̥�XE񏻈�e�A~}Y�?���qC�Թٰ���I�&��)tu�5h���O׾�6=�Zr����4d<��&����k�Eb%���9xn��E� �����H�<��z'�U��M>�_T�i���ʹ+L4/O���T�����L���A XI}\�j��i�9��L/!dG���6�K���2�u��c;�1?k�jQ��R������}�[��E0���Gd�+x��{�s�W��
,�����X�������V�y�j��ʵ�r5_��Z��6�j���;X���ȁg̦O��`2�h�ɘ�:�e%[r�ߗ( ��U2������D�N�F�D�0��}Z�,@���h�ya#��\�����,5m$ �)�%�efiq���y�ݸ�I��,����*&Y�C]���Q�1aZ9�~�S���{@BY*UFY�_*�Л�E��؛�Bs����}Vz��rf��P5/�@��TM���ۅ�voZߤ|��������$ ��x���ɼ
d.�2��&��h�/}�J��-�	�װmclK�Q"?�v"�3�cp P�;�Oޣ��B��O��5Oy?X)K)�5���P�@��qY������>E���&��*)e`J��e��2�l���}'4�\��x��#h�b׻|���6�����n�g�)~�8�Q������C<���j�Uyp��r�lx�Ӷ�kt�~�� $��Ҏ��1�a�g���=����;�L�@��z6Qf�}~��)�L(�q����@�h|��e���	����6�Ң����x��?��� �y�`��^ՙg�9KF�RsOq[�#�6Ol0a����pħ�z[9���D�"v[(�5��k)�:Ȁ���,E�#�'zq;/o*6O�2�m�֐�� �9�BÂ����P]gRF��	�>q\9l�j��@��@�e���L�Um �s����$�,��hW��|̘�E# ��1�<cS4�x�W^���ٹ5��nS�6LB���E�[߾X�n�I�M� �ȕ�Z�-�h1���R�M��?^@�*�\�_�@�Y%V��8rL��U���	�|�6�
�]l���h7���/~U�<��n�0�V�	�PM+8�C��z����	M�J}PWZ��Iwpgg������Zw�"����/���Ye�YBjW���F ��9cr�gQy�>��9�#KF�޴=B������Mz)+���V
�R/YZ���dt�RVr�2e^����Lin�6��+�1�iS��F�6��B����:����JWP������ �� c"#`�pÅQ����L͈Zd��_�2��d.O�"y��P`J��I���Bcm��!$^�ث&�B�g�CҞ%Aֆ$��d�� /��!vp�{�LcI�+���~����:!����¦��q��ث��;_�<�.�L[	Tg�?�zg�X�?�:b���l�7 ĵ��	���㫃�R�����Ό�8N�o�I�P�n�&�R���=f�~�L��7��0x���	�o�����XaH����䔯�:$AX����|z���`1|��D��MZ;�0��0�6GA�4�?���aߓ�GX��f6ez��dF�8���JB+~��@��T�
T���r28vHT+���yL
��*�'�����s�����!�?�\+u�:� ����m�xQN�+�ݯ�^�{��(ũb�$u��B'D�yε��zQ�f�fK���y��[ҵ�j 	��o��u�%����y�'S8h�'=.�s�F��:�]Kl��bkd�3\{����f)� �(fx#B�Aw��+�)^3�a�S�}�Ը+�l����}az�-��G-�[�2��8H!�ZE�ۑ�Z!uċ�߬Gn�K\؋�ྚw��r���TCQ�\As�������9��ԡ��h�x�>0�����5]`L�%1
����dN������6�=p��w�G0����L�d��L�'�N`�T
��0�X�i�j�Fd���Doh41z^��g m���?SW%�y����df��y�7��(��M����=S��R��U�n��V5�x��ܭ��="����/1�ܺ���R���>U�q�#<��{n<P�T��,e�:��T�֪�y�Z&~��Յȓ{���)�L3��=�R^���&UM�ҕ<R��6B�DV�M��{[h|N{��^u�[1Y����}�[��g�@��o����ګY��M�铏d.�b���ǿH�P�� g���?����Q�E��ZvdD4��^'z�(�g]��(��l�Bx�$9�v��}�p�]�`"�Ï"�@�N�T��2%L���z�Z,���l� �A��2�Pw�N�yw�!�0R����o�۽�Y�P&�'�K����`f��ƅ�j;���J�Ck��<�I�>S��&����I<��Ԓ}i��54�.M�ݸROdz�LҪ:��SqAJ0��/�lu`7ыEu���	b�8D ���Q-����3M@Q��0���J�헯�]"�����u��a����5����[,ˏ#h��k�'R�g���.)n�F1��D��L
3��j��y�V5	�Bq'�Z��0�k����x
z��B�d���g�so�;�J�\���k�A�z�JZɈ�oW�&��c�E d�>��O5��N���~34��@���P����*�`��R�%(�|����Es��Z�B!l��Pl�/��:�ev��y�`$7� �Ë������Hv!<K՛{���ϼ͇/~���ջ�bU����Tfe�[4vbE'[(��v�?\� �Je�u��עO\���,��s�+�R\،	�� �f�N0���f�Ч�8�e�׳��~�̀V�A�h��S�
X��jcO��a2���O)�fsV	5��T[%��'�3���|%z���t������� �r-���Ո�,53�?֓"�/����V�zD���.�~��5�s��וi� �TOt���K��S:�����m��M���n=���VRq�+�,.;��ĩ�߶|H�D�����9<X�D��p�X������ė�x1�&��ǻ$)����i���_� l��Y�m���,z�P��g�F��'�PQG�"��G��\�<ļ"�@�V���Q?ò2��l��$ ՚�/��μV���Ԅj�.%���C��F8APG��
�OQrf�./�0�Tfk3��Nɨ��2�ȶ�Ĕe�26 }K,��
A"�n���p;���>V�q��%��8�"z>`6�ϘD�S�y>��9B>��XY�<����G�gn��[fZ�$�ޚ��;���#��˭����ŉG��V�E&�����ͅ:k���Ɛ�!����;�g�D����+�����K��v�*��D�A�D(�	b�bH���ű�"4�ug�XQd��'<���"ޯߓ��˭��N���'��=�ᐚ�,^���YuC�g�����S�v��
'pY*C�Q�`�P�h�����@��̦��QW"��%|�^�/�[U(rV��Hn���k}�8�$�Z�Ůa0u��	6�2���SaǞ� �#,�dQ�Ƃ�� �F>�����v�o���b�q?<jB_d��Ĩۗv+0��{�_b��o��>���y��-߷�.��ݖ��5��#|;a�fV.�G8�D?�ʨ���Ph?��S�u������u��C68���`Q;����w���7���G�A���iÈ�7���b�g{��T���Y��K�"�G�w�+�I���ig��QW���~����>��+#�-� 9u|Z2g��,sP&ʝ#q5��f_T/����?�)�=9�I�j?vx׫��:W8j+�`M�����/lw��A,��ʴ�H�P���+�b�S�(�F����Ӈ���l�oA�eM��$xr�f|HT��2:H&Xx�O�Mٻ\x A��kʒʁ�J5���U������nR1\�m��}�+������H�Ս��jTuK:iч�&Qˈ�N�mՖ��e�n�5i^G�
�sO|oO�~=7_$A�o�H<-�L���6&(QA�a+��wF[ԅ�/���8��:�D��.��t}�$�u��#ΪS�#�#;���K�>.�#�kh����l��%����(�z��?"�Hw9B.��|�� �U����4s��ak�|��si��_Ҭ�f%AY�Zȴsd��z[��Vm�6�����2kp��e<�'	��eЫ�Ͳv�q?�{�Ծ��#=[�>�1�W,�k�2�^t�L뮫	;o��j�3��.��߮9���<��I�ˆ���'��c�	�i)@�DV-h����9E�1�LgU�A=1+Lj��)���+�3�C+�i��Oq�Oh�����2g��ОIF�1�ox��������ۦ>%�_�E�Դb	�U"
�y�e���Ֆ=���Opn��(��1����=���oa��E5�OdGgg����+���w�
��+|o�#e�hĚfi*�҃���;��8k)#��%Q�M��hG҃HH�f��ۆH�߷K=��վ(�k�?jcuC�A��{Z����|����\�yQ�m���L#�Nf�i��d��������ZۭU���ɔ�i�����Zx�Q��Vۍ��1��Y�D"��_QYzW_�������̠�;rV�e"n/�%D:�}+;G����Ub���$$���M����v�E[����O��FH����ZׄIg>+��LA�o��r�J�.8*�H�`׷17�x�S��63�i����/̯=�.=�^u�]�4��ƺ��+�k�nXҿ�ʍ�J̙�����l����F1k#�d���~ؽjޱ���c�۔gKkE7����]%��I��V�α��k����=+1~(BVʒ�����MF���O%�A���JRϰ�t��y,#R�r��r�Ev�%`E�k���7!܀����V�Ղ��:���&�
��S㎂�i�.�p*�t��g����m7���H����F�w.�:m�*
�{F�T%��Z֜�{.�SΞ�����tH�����Qd�vV���*����l��!x��;� ��^))k���F������"�V��u���g����	��E�q8���C�e��p)��}��E(��9�Տ�!�=���ᏻ�#�ɗs���E��4��5U��f�PK��&��G�i��:��5,��?ƺR��(-��T���Ty�g"�7��>L�6��il0y��*���Xyr0�2O���=<P�e'�&��'�2g��Ky}�rO|+P|Pf�� ��p�7���Tǧ�ޘ]J?S�ꨊ��;�s��2N0�s�)?UdU�R�2²�C9����um͌��Ҍ=�XЭ��X*I�7�h��A��Eh��)瘶8p��"���z.��G�W����㾏��~�{A["�զK�#F�<��t����=ꏷC̷���Y�.���125�_C��Y蒪�#Ʋ�+ʸ�� �w�.��{�5�2N�-��C?2d�z��j�?��w��|�c��]�0:t����nu�_$s(?��f'�X��ŋɪ���s�?���)"�BaӧK!���9N���z�j���<�3�3?&�|���w��ڜ��4��ˊ���������%N1/6��i;�6=�U5�$�ױ��g�B��mė���E��f���*�yX��&6�A�"{G� `A�����jE�$j�;�k�����M��ɵ�_I*�&�5�7������(��(-��|���8�w�����~P�̣���n�=S��:� ���+"޶�1���Q���C����	��$���>n���d��#�'"2E*T8*��~���㰥3��SX_��S�{Nʌ��츐�{�����ȗa���j!�r{� � y��'_�Z�*(��H�,,�禷Jfw.�e����K/W�|H|�
y?�ueG���d�J%Rݥ��:E���eY�V���ЩJ�vc�n�nų�hj��� ���Q��O����NEut#8f�P�S�WC	{QԔ���~��.Φ}q�ᾊ��$�f6ŵ=��%u���������6�9��3©lN�JR,����꜔v�7Ek� ��.:�F��m����(�%<�N��ëEÕ���tB�w�^�򦓆_�H�)gF�"��	�� ������ E R+�Oݩ\O ���M����
lP��d�����9.���FTr	�c-&�b�Q��!�j�����Z(5�������Y�Ca��Lw%�ްzx~�?|�8�_{qT���n�E����.������Rՙע6��wU����$J��㓱���_Кcvs�����������4��;���}�`���������{��zL{�_)�j։���]$[Q�	�A��#W��� �×:4N����]s�T����%*C�U�3�:Ml�n%N�l�k-#��6�>I����p���;j����Sq�Xr����A��?�[Խa',��J��A�W�o�x�*=����O÷NJp>����D�>r�IGҍj�9�
��H����0��n��ck�`�J�4��'�	:q�U��"�җ�B�D��)*p��֧d�&t�T�v,@��h�,�eݨ�Q��Z����a��Z�p����1�N�M2]mh�'3I���3��w���2-�t�7��cSW�}!	Ee�����E$u��uN10Q�1V���Tʓ�KYb�T�p{a3z�kW�2v����zs�^���˺�]m�󰲔S*���4���o��E�]�w���o��Z��Pz�ˀX�c(_gO����D� ��wj�#yX��d>H�b�˸Z�`ΊcYl�J�˯��� �//Z����M��h+���'����
�]������H�/;�K�?��uTsc�
l�����s;\�O����D���Am�-�Ͷ�>2Ą/Z��[ :vT����� 
7�"S+��cw�ʊ�Yr9XFe�A���إs!�����Qd�mK��v����Do�K�Q	 �*��ƹkR�"�fM�i�a�!������+SO�<�a5BNZ�	��^OE��zL{)�˹X�3��`��<��R��1�휱¾���r�����
�ϕH��eY�Amw����*�*�
��	��Ƽ���Ѱ큚�	�%]�O�m��XR1�J<::���z]��.
9bĎ(�:70���D`d9�U���Y��V펉��`�/!�X�Q"Υ!��P�yvqU�WD��U�Єk25�~��g
oE"��4	fj���r������ ����["���-�x����h҅;���F��-}7w#	SO︑�]O&+��0u�i�'��>�E�>_7�5,%���a��K� />��3>��������s�
�=)�/-��".t�.n�wo��P6��L�1�fR�۸�u)s֕u����Z���֮��l�H���8G}`�R���7p2=����v����Ԋ_-s"���X��&�I�lT����@�C��I��J�YV�3�����T��yO!���h0t�+��`�"�]��y��G�K`��� �q܁����<\s#J�r�z;#�fe�=z�X{���E+�8���M�����6F��f�S߈Lm��bf��=��Vq��Ԣ�~I/�|��MIv{7�!��k�f�F#o�8i��^P[��@�؆QR���[� �W�vI0<p���s�kӱh#��SԪ6�	�f6��V�a@��P+��e1_�[qE� ����c����I� ��6w���|/���^�|r��s.� �xoD�V���E�CI����YxL��:�F���)�t�]'�YǢ^���14J4�}�0���z�R��W�����(v1$Cn�$���]�p�pz��.D��_5���]I%����E���$R��p�4�yy=�xt\=�X�j�z�&u�2�������7��?9��4׀ۏ�C��9�E�d����-b6�J�b&����͂�s�v)�����F{	�X��;�q/=��7$V�r�Dtf��d�����`�q�#��>�.��Vg8Ç�S+���D��*K�BT�^ݟ�l��UGi�x D�#�%}np���P>���:�Q��`���"�����M��9���rv�?�7p���J"�o&�(x�y8r��d��f��^~G�$;��U�h�jz��N�3��iRUA��
dk��w`-t����\���{K�=W>��k�S�8�gD.�����h�w�ۮB���!���.���q�W���b��O�T�9��o������]��QF��@��ti�?��.΁
�S�6-����������3�$�Xg�!�{5<r�љ�X�Vu�h�2`])nS�a����dY��r<�:厍.��Ϊ�V�i|��oqhX� Q��Z���]o]��>��<I϶����ˊM2]��Sb���2t�u�䫵���W�Y5�8̚���h�I�����]h��O�3���55,S�/������M�����ݓ����w,=��v:�H�׺��n�@��[@Q	���#����*¾n�N>4mm�D��ڜF��FbH�X��=�%M�zd��W�z>S�l��
Tw̓i�snR�x��I�I�9U�0�t����V���͇����`�1U���JG�.e�����~���QE�%�H�s�O~ 8�9���o��\g���C^a`�b!�Yu��ȅ��X��}��P�!�h���펱V4���[*{ej�
�4Kܐ�TՃ�?�q�X7��e�������$�"�l���+�oS$إ�ڲ��GUGJ���"?j-�$��L�m�Rm^�fN���h��࠭[,�P_}kSfi���^7O�=��Ϲ!#����9�1��j�D��}�c�c�+�5��P7�S��b���zҼ��k��t\5]�by�`;��s�%�t��x�8�f
o��<�X�t��3J�}��[�rX������+mg;���0p0�4'��v2Xދ�;���ʩ!�|�� �>b;�[u@J�WwA�|���5�vd�Ea�K	�4�.�f�~M?�D�RK��=�Xjݷ��$��.�粫���/���O����y�B��W���G$���6��K��( @�� �IJ�o�xƾd�y<l��-2��H�2*i2 ��z-ʯ�o�c\=����t�jRǯ8�*�L�)�Y�#�0uC�S�s)j����a�U����b8c�Q��=x��i]�v�(��F�OG��X��J���z��N�z(+g��n�=�ڸ�K;����t�/I�۸�{J���y�ޜIK�p�2"�N���RT��m�����gN�&� ��C�7� ��������&`c�aDՐi���DBq`��?_4����4��ok���v$��=q�C�p,L�@X��o�ɨ�]��I��HV�E;}:s��'���v}��h��|����S��1M��e>fsY�iG�G4��&��/So�6WA��V�V��ꖐPr�-I��\:�/v�Y=�B��!�Z����>z�\�.g߂B{O�>�҆ �i+Dx<����B����0���W|����!8���1~�\$�ט;ZR�����ä�p�$�j���aI��9[h'�Z��o���|Z}9�oO�K�\�1��T�tWW�����n�E.���C��U{D�r�B��fqQ��H�.ʇ5��V��i��Fu�h�j]�"����ſ$���EDZ��]��#�
�(E��2�ʤʲ��u���>	6���l�G��j���X3+蕿9����v�"�6/��W V���@��[��s����-*���־C���o�L�g����Ym�`J}���0��"�l�
�P���W��V�@O��M��@��R%���:+���1}�����6���'o�0c�Y��1��q�ߟ)�nt�����gJ�a8�<���z����-��ui_&��A-����:��ѠW.g�\��Q-5)�^_&~�Hk��9�q_>:"�W����H?ϊ|n���d�\�>f.0.Gᡴ�r`��a�|av��ل;��'����}E�u����'��n+F@Md���X��;�Em���Q��-���<.��͘��N��ջSW��g�2���CBxȓ4&{Dߥ�PJ��:UZ�p#�ѿ�_�Z���iCkV�ayH��i��痪�����26Z�[�Z���?A�R� d��I�����*�R�Α�%�Nĵ�ذ(���R�&�Q�B�.@H�=O�R�J�J2I[�m���4vF�'Ǝ�k�R3*x�'':j[C��w���u��g�`�\Y�Bp��N�������EY����p��N���V��}Л�����t5�9��k�#�}�����p��_�X�/���M�x�E�!�曥(7z�]�3��2��epUr�%VƆ]T��rnѾ�=4�GP_xJ��t�L�������3���4d�>����;�TK�/&]<�=Vv����Nf�S�<��{A�W7��p�'��?/�O�et�����7����n�L��10���v��H�0]�+�6�u�>��� Od\�b�� �U��[q���g\V�ۧr�˘�FI5���֍��v,+��p3�����_v%�Xx�x�j0h���]̏�c��N�
7��8C!�����lr�O�r\��,m�h�21E�2~��~1���`�iyc�p�a�*Έ
������W�L<i�Y-�8�ƈ��q���v�e�+ i�Z���k	�Z�L?�o�P��fՑ-X�Џ�RsKdFk:pHH&�a=tq�Qtw�Z�6�i�Ԑ"�`q�0TN�Ӻ��p(џ�����]��g��u:拝NԾR�����c�\��f�S|�>�z�*��ve.��_y�2B ~S�9�3(C:�^�����eA����4��C����+�+�$�7i�R��M�P���x��%"�K�$?�(���=�@#!�b<�S��Áu&9幄	�_2Ce�2����w�{�>@y���N|������cV;!0n�[u-��:�x,����@�^#S��[��`�'n�H��J�e5�� P�����\��?�"Ȝ|�w��=��~@��+����K��}z���m��i�L���["�Я���x�r�Y�S��岯�x���R4����ǚ���џD��(l�r��8 M���ʦ�!=9�j�/�,F�c�Z�|���H��U	�����ھv<O��W�f�,)ݳ��C@�edǷ3�F�u.|�r�M"9|m�3���z�)�3�e[�!Þ��(��s�wL`��I���V��3��� ����[z�~�A���%�MC�1����R�0�������h'b3�7�Z�.��'���0��ɬ��Q��PzvZ�m/���:ޑ��t��k�׌�/:K��5��1��Re\e ��^�_6N�l��F��!�+Nk��Fh�G�{�'1����?E�~�I`=������wK�k�2Z�=J��>:�Ģ�T���˩���l|CkD��5���	W���.p�N\SY�;����<dl\..�b�/�i�C���<��8�����T�{�k��ws� >0�W�P_	"��˼Ź�9�?V_7����q���i�#�O~�^9�JV��XTϒ\
0�QYl$[hC�>s��ŷf'b7>�P��Ӳ�
f2
��L����Hʁ�������.埝��}�db�l��i�pϷ��w��W���lcb���A�]���5�����0�����z���y���Q��U���.��'J�@E]-��;�Uigm��x8ӡ�1�� OᦲJq��� �6{��\����8h���vX����H��ݪ���rgy+3K/`�/n�����z�Ԑ����&5X�
���o�H����=W�����6e�����Cl|��P5��e��'��AI�>���8u�~ߦ>�l�Vj�%��2��Xa�E�����%�\[6��l�4�{����0"����)�e(܄��5K����M *o�ߠ_K��׏�h���+Q5�<'l�P$AYH�}J�vU<>x�PF��=�.��,� ��Qy�s	H����o�d�Hn���l�l�c��خ�}��{TcB�����>�1>z�e�0�k!ɨc,�p��b���tK@u�Rg�8���@�;�<;ѿ]���ù�a<���[<iԙ(�1Ddg�3F�H� p��̠��9��D/���Dewr�ZY9`��V��>��Em2�6��v�ڀi�y�����?,ç+�yX�^��`���$�|�m�r8"�^����u_��t�(�L��{��R�њT�o#'�`�6��ܪ�L�FC �7�w*�A���y�h	�wa�$]=_���G|:��f�͂E���;s�ء�R3P^t�Xw�����?�����>���lυ�TY�%l�S����3=���q�K�:��+	S�'3�����o2�~�z
��69�*��!D�f��� �lm��?�|�/������}0��|J��RR�F-��D"�4���WT`���B;� V�����`�����hM���2�� �z�܎�N��qooR���{��^���9��ߍå6�(΀�� 2��񘖢1�M��	��7e���oI)�Ǎo6�]��n�JI�������ޚ���[�3~�ʸ:ks|ܾ�j����72PS���q�A��0	M��*��1�r�f��|$�� ��QS������|��
0C��Y��:���_�霳��N���&DJ���a���]w)hC&�$��y�rx��嵐e�j�,�-��N��<=��u�k0(�@��p��9��v�v�����6���BR�!�=��7��C�"�(e	`��<p!���[�H�Hi�|�������B:���/�+t�����83I���&�A��k4����v��P BG1������������;?{������%K\�Z��I�Ѳo+��8ybwg��zt��V�b7���y��s��ˬ_[*9?�)�xr��m���R�0���XQͤ=��gJ���mgXS���<s�r+מ�ć}x8;����wF�W9�f���\����!��Ᵹ�.�𞞳��C���ю�k�I��	\�����ߋ�������0����w�Tt�k���x!-���Ɛ��Z�C3T��˱���.���*8��#D ��R��1p}�vӑ���T�s �]z�[-r�&eƟ#fe\�o���bj{���>��QʯC�e+�ö_��fy�s�h��'|Bb������_�C��nY��q�y��`D�ӽq55�"�&4*_�/�}����3/t�dJ3����	��i.
�۴Eo˲9�-��� �M.�����roG@�Q1q��Mb�KDO��A_�4�9=��3��v����i��; .��E�� ����8��`�q*t�(V&��8�<�et����u]�.�7 [�:��^J��X ��9Tz�V���k@�
��� �Z��}��ymף��~�_��^ �r4\l�����O��5�xVl==0��jyN<8Fp�l�!>;#ˉ�mװ�1�h�5�8R?�J�MW�����w��2�j����hj��޴X,/
�p���H��*��'L?��j[)�2(�.|́]<럇V_�_���X���Fx<qar������o��Z�1U����!%;F�"U���x�ة��G�[�lH�������%'|�T�u0He����P�|H�4a�d=-YP�7Lúa�e��$�� ~���^���KZ��g��Edu�)g��gS2��)�ּ<�����	]�>�$8�O��=���7} �{��
lI���f���v���[�!¿��q�v�k>�����7�SSқ8����hC����c@BeNS�x>�ޮ��&}P�e��|��ư�L&Q�2y�m$oTu3�R���탃[R�(F%���}�S�乼q#)3I� ��P��$#%�)���R�Kp��ƳKx�#>X����;�}���bi_��+C*!'�!���������01���{wO�}f��34h�;���I���-��G\�vS]�Ih�2�ߩ�_�YR,v�o�� ��ᯔ�{�Z��ο󁎉[xĆj���!8p��M�_���ߋ�h������j�7w���PoWI�I\���p�@Q�،�x���gk�}���������RQ�J���q�)�qz��Z�Vv�d�8�$�(.H9*�>����7�͝\�j`�To��l3�����V�SW�o��D�Y��`Hܑ���>J
���hp��a3N>�NKc�� �w>���J|Z7�|�ZS����-)�a �,r�I��.a�+U���m�+�1��=o��js)o,#ٕ������'-r]�W2���lc�SU��J�-���Iߙ����3M��B�֨"(��έ��ŭfl���T�� p}�$���4-"ÔR�2�Ѥ'�}7~]��Xw2��FB%.ڌA+L��$�7�
��#jiO�%�Ɲjj�5�!�EÕ4�N�D	�&<�\v�+�1�wr��&��ID$G�ǖ�!s�S�[,oƝ��?	-g_(EA♯���C���dKl�]6)��w�hk�IfX�����%i$�G�|ɍC�W$�0�U˩o������A�\�M0p-%�U��i;��d�K�6������H��bhK#�A��ً�r�e��9�:TIN���G�Kj��
4vɕG�<4��"J�ң�8�: ��TV����W%Jk�
]�K�,%ֹUj�+�U�p�<$�R� E������ �s®:$�@Ҍ5���~*�Mt���&i�3b.-�WNGE$s�r�bN�J�8s��NV菟�~<]N�z��)0��r>\8����_^G�!�p]��!���Y���>c�O4�t�<5(��Ee���j���ƇM�ĢmlV�G�!5%~tj�H�Y�C�
�ý�>pP���pϖw�+%��_'�ؼI��Y�D��I�����"�'��Ә�9Y0�$V�zZ�Ӻ��T,hZ+�"�~��hL;�SsH�-{s��m'�S�Yf�V��P�Q�8V���:��mR�j��N~�M�Bs��Ј��]���v���kh���*51*�S���خ\~�G���A����Z��plI�:�E��lu�8;uβdp�l"v�B/�V@��q���/��7�ۉvү{N~m����Qeވp��t
-���@k�i
�w��:+�#�&a��´'j�O�{G�p�Đz���/�^������4�3��.t���V�� ��I@�p�`������=eX�	�ۚ����'�̀f��/���,ީ	����h8���R�R�P��kd�fx'l�l[ڜ��D[������bQmͅP�27�u5�k?������J5�X|x���U�`Ps�d��+]��t�����VI��ۓ����@���],���)<ߴؓ_�H��@O���
e**�L	�δg�LX�3��ɾj保e /�8zaքϮ�8�Qɒ�k���>6A��~3�qM`A ]_�K��݆�,�w�_�=Q{�x����h4q:j2}�߶��9 -���i���"dL��;��P� �E�/�bI�x'L�8��M(�0���k�G5Vu���G�7_Dw���>~Kc�,݉�+���DQL�b<�� }����A����e�@�Re
�T����kO��/(p�%�b�+��C��`x��.�LDP�+����t�tl���n�1�=RΜ~sQ;-?	kq% }D;^�I�.X��C��T�ٛ��DfYy����W@*��񘕕;�[���(�F�df�8��M1���Jks�F����U��&�<3�ƦIK~"��,		y�R .H�WBP D�W���q| �4��/�(�����&QI��ÂYY{fl��3O��N�G���B���B%��ؔe�ڱ�t�$SR�>�^�Ǝ���*Ϩ����J�COh�$�0���0�+X�L.@j&j>�z	6�"��8s�^[�&�3����]͋i����ۊ�:�F)�1] �t��^
/��RX��Y��|�8{�(8�����z>	q����� ����T�? �5v�R�I��ZU�Бc\�Pq����_�e��
/�	�o P:T��dT`OU�-�{��Do��b3�B_Ț���iIV;7n�N)���g@&.�5��"<|2�=y�a��^A�̣�`�d�}�%���%\#y���yث��P�õ��Mk��'B3�0�r���/���<d�^�D��6h��9Η{�|�۱܌Yy�;s���z	���cv'F��}m6�h?�����Z���v�kP�y�<n����s^�N�dfM�H�}A�H�c��lRT03�]$x�ψ��F���8�]3&�0���K0,��Y�/�J^߼>I�)����̖�S��X��>��|S'�����!bے�ťe�`�>!�~��~�J\�F�p�n�بaB%�g�����Z��,U�+x��!�i��L��4�!x]��!��4zO�(�pɴ��׽���e�x�����0�⽶*"�?��|�����Z�I��o2��=Lˉ���������#N�t���I�XE�p����$%\�|�>����-7TL���I�5(�H��(�k��Z���ֱNα��/�|��2

]v;�N~�3�mהj��@�>��Tw��ёt8�U�/�B���ٿ���Z��FX3�h���&��7�g�4r�9z� YV:�ӊO�&Ųr6&ӻ��A��|:q�,����"�ڄ!O�؁i�>'K>�:p�C:�O��P�<�n:�V�9�sh4-��
�㹈�1�lշ��u�W���04i%�"{����A	�r��)u���{�u
�8 �Cс�ɡ0�I��E��@G<oP��M���a�)���'���Ar)za���H��+ǲ�
S��A�gY4��p��	oU vS���Ne�#��e+b�n�/��U�D͋�!n�����k�R��_��R� 7_�om�S��k�F
�>>��E������4:~�H�t�J��L8278�dkh�8S���n<�)Q��Mr��b2����ux�/�b�oS�4����D�eU��q1 M�̕e�q��c��sQ��?���7�{r�l� |�;熇�_����ڵN�:|N�O��H�[K62�!3���}S��=O�C���n8\],�L.]#G��~u��G�˒0�:��(|:p�ݡ�E��J̆R-�̻(�7ȝkw����oN)�qF�C"])x��	��^�]���U�d '�w��t��b>\m�.�8M�HIvЂ7k���>�����8}�#r�q@ZTL���#^��k� �G�/�9S������W�c���ar������Q�ry%���^!��?�e�錔7���+rߍQAH�Xp�iΦ��i�3�'�� ����]}O-D$���n�ɻ�%�`�d2r�YIB� ��=�������\Mv��z_wD~4QUr�N���XL� �X,��<�50�pf|�x ԜE�G�U�Ii�xH?�q�>`�K�)-��е��KM9�?��cr��-W{��e-���G��¾���B/�(�[�L)��	A�I�||.�)ڬ$���ϚgR�qY�v��=� .��sJ,K��Y@ܹ�n/.���FF�yC������
���h��h4J��M�h�ј��"-���6TR�Ն!5�~֤��pTG��b��"G����J$����zp�EC�R����!������(2]J����Nnt^h���?=IN"��Vj����U�D֐'��C~|B��f4+�����T����4�6��~���c���z���1�����񐅮	��8cB�����������xz�2�M�G��
�)����5ÒUKF����]���G���3��B��;0?�( ���2�P.G���3h����v<
؇��}����A7��Wv��XJȝM�$U�7V��~PA�C9h�M��DͶ�@��	t�X�NsB@	L{H����[0Iq� h�`���k����D�t���T?��vUi=���1y�D���������ƿ1SW�:���G�לV�D=���x� �� � ��<��'�����F��;�[���$4������~�>qd"����.�2��%��R(K-��#Yˢ�E)'���:Ǹ���d.za��S� �i4��Q�ٻ���� �~t�M�I�5Oj,�Z�J�X�@�g�s���[V��}��Lo%cC�b��$��^�a��L�cM�Q�Zl$��E���=�1=#���ć���6A�!s����K�l��n���Uۋz�ҚR��D�PY�QI�Fj��|��t%�y����pI ���X����r�����r���=1�ʭ��ί�Ăw͉<�) ,gw+���k�P��r>y�4U����'���'Q���JL������l���'�� i���#�a7��N� {��Qk���@�E�TLm6P��j����Ѐk���a���I���j�����Cg�u��E	l������w��g�~���F>Y��h����q�S��z�0<���������%N��!'EO%e�$�]��O��Db#����:W��/Ψ�90�̀I��rf���}��C	��^S��d�q��C����.�4�����L��b���ڢJ}����c�-3��Չ��~ ?:����g=��[mW*��quI���N���7]�r�~`{��Ƹ�{V��l�J��;~�W~v,�u~CQs��i@���˚��KEw=rɁ^����u��Y�4��09-h��c��'��a:p��o	��<,�>�כ�4u��'~�4�l+�7V�a����I)��l��
�͟�ic��t�h��9>s*<�:� h�J|�B����!����Ev�Nz:"Y���ٶ[?vet�㋓��RSMs�g�9:!���i�@�<,��� {��:&�q� &�c��:C3�o^�k)�܂�M�=)1o����#a�'ӄx �iR�\�~�̽��T�B%�2,!R�/[�?�<�dC���K����#Ъ&@�$��N$j� �)s��o�Nrq&��T��>&o����O~始��[|���-���Gu��U�W�̵� =��~��i_f�NE*���r�}�zX-��d��k>",��\��χ��K�����䮒��$�q���C��	Y��䱒ev��)�e a燶��B�]��h�Q���o�c0�
�S�]��B�����)�������KȻ$q�r:�q�6�t�,j���8/�sa!�2Y`�f���\^ �Į.�P蓞O� ������wGe���D��XS�jQ�c-��!�� ��|/l��l�>���i������,�r�Ȱ�'�{p�gH{�#���h��k�}���C�4i&���+�rq=�1�;^~�]� ���B�� �dF9D@��1<��9לfn¥5�i-0ش�&4�,�4�/��.����^������
�7$�^xO�M3���!/E��CM�sv��&V�iTTP?�4�5�RpḂ���
9��zw�)P�p�w��*�s��#@PNZa��
��#p�����P��F�d}��0�tH;�q(k?�����= �3J�Wd��Fj�﻾>��"�zRJ�q�@����dMɋ�� �!��	�#��o�A���(jx�\��e�DB�-37��z.�i�j꩞p�����S~��p��cy0g�Nw��3��k�_�f�ʒ<�(����w$��J�9_b _�ʂU��)�f\��M0%.�l��~j���NKp�B�"�4�*|q�r�@�C,�Pz��Nn|d��؁�����9
��
�tLǴ_�E־|iZV��U���NƷf!�P�p��5/��֟pM1L"}�	�`,?�T�Bj�;�Ņ�[S�Y�n���3�i�D����0�W�P�{���4̧�^����0k%|��U�BU!2_�&w�-!���8?����G��m��yO߇Y��V�S[\d�5�������=5иe�l}��� Lq3�j��������1?FW.��R�8��}�X��\�@�����U�M@O��M4���%�yk���Q(��cKz��7 ��P��ݶr_:�Ս�{������
}��1�1�Sq݋M�j���.�� [\+0�Z �be�ȼ��W'_�vTl��PrPD��Z\�U��0��wz��W�ߙ���B5�.. CmZRַTkȠ�9E�{T��@�;47Tc[w�)�@;f�x�E\�F{��y�-f�I�+s��M�Ua�
%Z��'��ɒRyz��1����;&FS�(-�/�	�J���8b[��Km�>Ǘ�¢]��0h�>q��l��4��s�zQ_P�b���q�r�s$�B�0x�B�U2}�8��c�"�ɺ9�ɚ�v3�L�t@�5U�p���R���hY�g��o6:�#f̋�e���0�,JP*đJ���E�D%���\MAbgI!c�)��L���o�:�4z�(Y3�d\��v~Wĩ�6"v�H�� �qh�"�y&N�B����H��Z������_�F�󞢤��%� �4�O�$^]n�%�c���t��	��7DĲ��`'$Y+�=3����І�������0�:�~1����uui��4O �B��f�씒��y�<��.��qʱD#_l�@�=��Nb�{9y��\�R�U��eX�h��o�b��ۇ@"(���s3Ss��GX"���|���^���1i��}o��JAl�C������H2�?�����D{�ȋ\�����g"��rL�Do� �S��1j&�\ߵԭ@�����҄��Q�9Q�=r�ggz׃"G&^X��Xc�M���ű�*�ߣ��tc�b��UKקIw^N�3_��Z�+�uk����E�V��y�.������I˛��~�^Vs6�X�Ed��m:�Oj�_%jˬfP�ßp�Wv��>/g���� 1�-k����j)'�6�
�>�q�ݮ�ߐ�a�P�~c;)�H���)1黄`.'X��nzy���<�v>��2�3��wMO߶3?��D��m%�jl+v�+����N��]����'@�����S1ۯՇ�G��͡l��(�95�
*w�$�~qhޞ�y�]��jx��{+m�yq+��Ƚ�;�#�G�K���b�a�r�T�p���
$�� ���4��#S��U��e�]\�!7���|}�rg*�P|Cs)�+wǇ���w�&.�v >~	gg hex��[���eɩ����h�|�Y|��qBw^@�K0���Q��3�Ię(%A��w���_,s�Le����q2.E�K���=VJ�X[ݑ�̉)��0NxAI̟"GI*v�쬶Qv��2+6�d���>�?�2�rV�e�1>qBZ��^�r��%J�����6����1ٚc�	���;B|8����A�
6�jt�5�%�4h�{�O3]��c�\L������٩�l�#!�r��VP��f�<
l�ĳ�SVW��H^��QxM����2'J��bCRw�P,~9�c�a�c	j,���z�>������W-�T���:c%C��;�2t��b>��O��gb_�
�o^yVY�����2!d�S��^���D0x�7P(�W?I�J"�I���������9Z��]�����Tv>�H��:;�ZI��J2AP�s� �I�#4��[E8?܍G�.�f����z9f0�gH�T��Ml=��̯ghL�=�$���t��0���������Q�(n��%�Ȭ��N��u�Y�F�꘻8�I�R[4��͍y K6��ٝ�i�^
�{������eT����+K��E���N�HDb�<#	G'��_�u=Ĥ���\�ڡ�;a��@�{)E��^�$J߽�k�ēl��nlf�5�)��o�O���B�����K����+zhq�BՅ����^T>'N):ML�_��z��U� f�¦���<����GJ��%{����xX����b������������[��"u��@�^����;wdH���e��B17�J��}��w�s�YN�:�H��>�ϳ�>�MU�-���N���h�ŧ��������9J���n�l�?~�cV�C��]#�!�&(����YT<d�v�.9D*R�0�Q$\C)���؄,ƌ2�
�sPYs{?�:�||m$O1z�P����8j��o̒ ���x?��c�^�>:��g_��ɳ�c<��jz��ѵ:؊��n������| ����
�"½Nw���8�FO8��%����*�1c�fi�
�-�o��9���Y�}5>�hm�E���n�����z�x�p���<P�� 4~g ��Ċ��j��}{����5Q��$E�w/;_D�����c�E�/��ߕZ:ը��"�=4A�i��#�}�3@�kےz�[${?��׬�L|�u�>�c��R=Yc�n�����QBP&�n´���B�t�;�'�$p���'���f�}Z�,^��6��聇�i���v8��	�؁���1qh�E�U��z�7J�M��|�"S�?E���}�^���6��!�K�t��|��D�鎲�~���z�ԙ/g��ڗWsTL�&`��$����a�x~&�LnMPwB�5�=9�`H9E(�0��%��B��ti�[���Sp�j�1j��M�Ozq������>+V)��T�LG{$
���IƖQl��C�ӴP������d�Q�П��]�J�ܘ�kcA0p�=!�;�6�w"���9R\�]� ���ͪ��BF?`�5QW�'��+4�b��"͜�[��g�����d���p���o�P��e����냿$�AW}"R����2,���(W�ƻ�8#���+<g(�cc�p�b4��*���R@�`x���Z���%~4���R��b�LF��Jb-ߋ�a��@������d�N�D�2��5�uw"�.����>v��P�;:á�[ni��8���2���벊��o��S��jD�7�wv�'s!*(�޳4�^��m�S"�҉��A���-m�<�7x!~�B�J9!X�W��ݣUo\$<�ܣ�Hd&�9:��^�� �����p�,+/y����إ?B����7m*�y���pN=�u�,���{�d�E��W`:s���:�C�K����yO`τM�gۋb�e�m�7�1|���9ln����YBR�/��m�i�{C{����5eQ�ٸ��\<�P��fh\[�}"�1Bu;|��Zr�R�Î5�P���+��b&�ye=��9��v<^���)��e�lG�ԑ';��n<(�!]�.c.�R��D�]⺝�|�<e��Y�>%6���U�S�&}?��t��̔TS��� fl�Q�`5�kp
� t�$Ku����mbI���E�n���%R�vپ\2)yz6�r�[I��� I��pByiY��1?�<���]�0�F�ä�}�{�=B71�������vBvgv�k�'a�q���������l�1�5,�hwe�];�̯ԷY��)�m�+V�o�9�qFzgM��r@f7x�]��ս��Y�m�����zQO~���ذV���:�����T������v��rk�W��q%cc/l�/�/�,�Ĉ��*Ƽ3^���t��WJLC� ��c˹���ٶ�ON�2G����3_�FF}l=�6:p81�;�y]�^2:m������a�h!����F����w�,��8�tʳ�;�.?<����Iw����nN}P8tǕ�x�UO�(t��;�5^�ڹ�`�B�t���dz�B'���@�Z1	w��VΖX�ki���!������w,U(񫩞Ѕ���|�][�v���pٙ����P9gn��![`�냦�?[� 跫ͩp+�8?�,����IJ[�-�$���ŔN���Þ1�i��6٭����G����2�8G���uK���&�����%[m&�ڔ�(�4�)�F�r���gc��9'�̝�:ɪ׭�גuӃV����7-�j�1��V�������y@׫��MQ�ʇ+�K�Ƶg��� ���qvw�x!�i�Qwg#�X�w>	7���~<֝�;��a,���c�e�b��1^�~C���7M�Iʵ|���n��u�P�W"g���A6~��]��vi��bu��)��-1*��9,�)���M���C"��l�nV_-�<�tܟ������dn���y�<K���,L������m�p�������E���"!�9Xi���yq���=�lS�h+3۝�l7�T����Z�v.��I+�/����)T4��C��9t�`��\o_ۼr�<s��h�޹��'f�@,�׎��|�#o�G��@��J��X�f����vx-j�Gh�\��4j�%TCDڧ�wd�^���T�Js;"����*C�����������m��+�@p�����YrG9x6m �-pF�|����LWԭZɫB�d)}�_��Nqt(�?��R�� �=i$[���`w̬�{�':�K��z�Y��+�'����i����t���A%�r*�����_�b4�OX����{�n��,�(�v�k�
�ŋxU��
�A�n�}�]F98��"���M��� �25U�`�),�ex�jC9Kj!�M����泑�?�+(D�޼=\_�-[w����7��*���E������7j�Ča�Q�n �YXi���߰-!4(��|<��UA��0N|v��KS��f�����>N.^i!��'�
����9-M3Fx��\��!1����j�1Ԕ�o���g� 4eI���h '���~'��勒������u ����'���Էߣͩ2c�w���u�r���Q�u���Nؾn/�
�!I� ��۵	!G7�gnT|�?�S���bef(Uh4�����Y�