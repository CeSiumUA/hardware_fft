'timescale 10ns/100ps
module testbench;

reg clk;

initial begin
    clk = 0;
    
end