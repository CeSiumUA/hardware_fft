��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�
/�Ast+�t����h��'��2�C�P����d��K(t��F��2����(3󜑽�-L�_�6S���c�;i�L���P�0 m��2��x濚L��EM(����im+��_t�p�A��ѵ�ȍ~���s����.[m�r~��:|NȨSм�n�.7�[_��h�C��;n�b݌�����i'�|OvV�/��ÑӐWCD�ʅ�|�ޔ�Q��~M�]���	17Gwu�;�Q��q���E5V��Qr%u���ݥ��^�9P� ~m�N����5���񆓚:�\�[}�2.w8�oB��}�O�]����e��»�z��D56m��9W��~��&	SSb�ӯ��9>$�����*?��a����:�ƹ1G����{����۵|�:��	��jo ��ir��ie��L�ya�{e�6�����}���¦���5����P�R{Uap��ɽq��<AxYf�_�j�P�aq��(Q��iaGzʅ\}��}@�%:���Y��{p�wҞ1��2� Y�&��Ī�lG��,���iSL��s_��J��H�g��0��X��@KR�B����ã%E���Ki\���M[&��6<�Ėk@�������kP��Tj��["v*�ķ��`tD ��}KًX����Dt�AU�Ȃw�����_�|D���@yXwx�W�|��+�Xz�	&"���k�����g!?�j6	E��o�c>Rmx:��E��N�vV���O�1;9�<,�(���2�sA��oQ�qNb�j�R�e���۠������k�w���E@��>�J��d�G���#E!�Bf�i^1�:KN�;�{��%f������[X�������=(XW �`�1��4�0�J7��c���[�է�0Z_�廬��>��x#�8�;w_Q0�|�7�_ 9�mX�@!b17���x��U�58~�V`��_6����\ݔ�rm��g���%d��:�"؆�{�l�˺�w�����^���ƍ���8q�xOp-��
S����-&\c�G[��&y~�kW�c�������p���Ŗ����k0Ƭ*��ӏ�*3�|��XK�O�/�M;�)S����-�wG�����0��I8qʆ�������K;*�A�=������;^�[���uxlw/��\�����B+�	����+�'+�J�+k�����n�>��n�ݡg5�`?P����l}� �|k�"�J���ݰq&����l�3\{W�^��]X�-p�kQc��F�OXZڒ�W'�"�/Fj�G��_[A<5�~z����b15���1K%��W�Z������O��^��?F�<y.�2 �d-9U������S�̥�������]!ɔG9aڒG��2T��]�zN�D2ի!3l��`��78;3���V��̸�&�S� $�R5��V��5����'6z>f"��bQ���omZ/�ң�m]��E,�
�͝�ũ�����]Z�6�C�gc�rw��"���bWDl��M�ʲ+c�+]�Q � ���q	��j�� �Y�ׅ�f��]W��@�8̄鎵;u��:>įſ}q�J��φ�`$������	E�Z-ܩ���Z���=*>�&�����Fm`N����W,���	c;����r%Q1�r�f���'�5�?������*<�l�K�`.�=)�;���4Ǫ�K�#ѥ��dw�m�̎	҈�Lf�z���_���@�n����P��HCjz��u��G�@���:��f�w�y])��Τ��[ܔ��{�o
�i�0���	���q�+?v�u<�����z
^�'�q�QO���.|}�o���m5�9U!7�@T*d�C�H&�����E�벀O�hS�,gV�`)�7k��۾����PBb�a,�}�fq����"���랷��f�>f+�Լw���)[ҋ؇(�S��Ę�zA��4&`y���z�4)�W^Nd�ad�����&���Q�Z��>>��T}��< l):�j�U�IT|u��Պ0�\��RI�ϝ>�eKN9O�8�?=�	��:�����ܢ�&����ۻy�
��\��7�j���w���������~+墄��4�2<�=���!��Ô[U�6��Wu(	���ks��&�|�uOY����~�j{3𷔴������ð���'��El�iljD#٧�\xe9�T"����[0r�.7���;vң6?���@!lA7�3��Gz�u;�*ٛ�������Z:zeFv]̰�zk�"��m�{ϾG�qG:�x.�R����96��3o������N�a�`XYp�9'��r�����͡k~Z��Q�d�rTB���{�Y�v�p��O���<B.��?LKQp�'�����I��㊺������%v
�qn`߃E�����ʏʇ;*��M����"��Gp���|���DC:̔6Za:�]%lS���l�����Or|�[�Ѣ���)�{����Dý�(�A�RnY)<8�h����(A�v��]���G�N�E��` @�g!�g"�O�8z���z�|��h����ЏW�*ؔV���ܹ�|�8��L�جyQS�莽�=S���tK?�v�����E���{똷�X��j�,KY�n�{ʐ����'�k��_�~��^��$l���?v;�
�~����7�?[�fAK6�Ǡ.ދw6����1�S���P���tٟ]�u9{0�p}��~3	@yl0M}Q� X�z׶�"�D���rO�S��¹歅���ȄAw�,&L�)B"���+zx{}�yF�+Ψ�<<Y>�J�\�K�"6�����;y�j�3��YQQ����a�+aCc4'].�po6�������6F�݈b(y�! ^�c�+/(���G��K^(D��eS�k�����!�W/BZ ����V�B��"�A$����/��e�m���e�Y95'0��3�a�ld���� �tr���W���}���I?'�R�;�rp�pR�.>2��aſ����e�`vy�=���vx�d���z ��ȶ쬮���<j����%e��2$V���T6��n.���n��y�����tȫ[\���O'���8F�)z�/��n�z�(��玀�Q^IA�ƪY5BR6�!3�M���M�4\91&bS�}�K�{*�����������^7C[�sYE�{�.IUN|��ǰ�ܭ#ìW��:H���8��-��!����H��������h���LtD����_`�X��w �O*�Q	�����?L%޲S;_�q��(Z�^G���=t���������VK��!y�^�h�a��QW���V�#Jw�&�"��|��Ւ.�&M�,ߓ���}��}�Y-�'������f�?vaw4wz����-v	7-s�@��вl�=�i�jԭ��#�&�h�(-� ����M�-���j�9�~��Β� Z�ˈ�z ��_.��-�y���Jat�I�9�kbD���t)}:���� �@����3h/2��<	"��9��=ģ���d�����?�k�^b�X{�L�s2(��9�"㑸��ur3�}E�> ��}�}Us{�p��D�4�p���8��$�Ǫ���ɭqr���Q�U��GL�7�E���	4�Og&{O�t��>�%P̣Q���i�{�ގ�$�^�A<��0g�=��:c ^��59/�h�V��7?9�hlp�*�N��wK��Q �S����}ąE�Ȫ\� >Ή1$��A0���'���k�Zf�=�摋��I8Ӹƅ��Z�B�/�\o[�P&�F�cf�9�de���,���,���N��T�q�q�G�'�0d"d{M��n�;S�]�w%��bC��0H�H��ֹ?��M��"�owO��n��n��\Lg>�3�V����#C��9�FC߶���)ͱ~�ȋ�u���,�=���
�+���&ڷ܎$U�7I��ân�IYZ6�S��� ��eﱺ;��x��]1ߕ%-ۑ߽�'-�o~C$?�HܻCc�O�^M�8Y*�����9ʠ�#60�2H�U�k	�3���8Y��l�����W��y��E��Hx92�H!l����<=� ^ϣ������f�r�Γ^V��?� ~;�"jM�z�~�	tE��fؙtHB�Q�[ۏ9��^��� )����b>�K�EY�iP$r�C��˲~t4e�b��+V��z�q�$�rf�����Pgº���C4ZȢ�	�Z��h/��A\St��A�-�;�l�N�^L������@��u�T�؎���y���l�K��;2��%�_�I0���H�� �e^:��6FCl�fX���sdi2��������0��ւ���0|^�vX�ػ,V2�Ge=-K�I�y�'am�V#��g��E]��YU�Æ�J�ۜJ-A��UҎ���B@bU,"����	r���DWcڮXo�dSZ����nw��v�P��ll{��,b��?������+Ŝ80?���&���^JZ�	�p�q]��	�j�z��V���d*X32�W�9vR���<=��`�H<#fӨZ�^�l��~qib(��S�2�F<�L �񭿐����0�U�*�[��?���dH�͕+.��[��s��9ǹ�W�)<4)�e���»�N_.��^=S������e� ` ��=%1��F� �w�R=a��������uhȃ=֓D�)�����e�]�iw(�і}O�-�����1RWV�֭�ʸ`q7	j��B=%����tk��$��TF�c/��)}ጮX��L�q��:��ښ��v�6���[�Q��8	�Oi���P�.A^N��S�dѐAp7a�F����!z�x�?��c���"�ْ�� Y�bolq|:��
�pqԴXg��N�a:MϏ83��rf���;:y�F���W�-<&��sh�������X�=J�@8�4šԸ��(li(�Z�ο�ݦޗ���A�9���#@
��4�9��yN_$�B��
�L	�U?q3j���������)��E�����A��b���'�1� �=ÆZ�ᯋH%�IDJ���[	��-�ʍ�4Ԝ9�'X��z���� ��̥������A���ZsS�{{_J����d�����wt��뚽�#���Jt&�m������P��b�W���Ԙ���Jh�,���>����^ ��Ce0��&�T��r�L�����z	}�SBi�)i��PЈI���C�[�L5K��.p���F�KC|��iC��]�qe�