��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�ij��(�������̫�s���֊v�@���PRĎ�cj���3�Ŗ����i@�y�Yמ^���(:~�]�%]��u{����jA�
x��[�}�1W���)�e���`OI6��bDs��x��`؜c�Ǘ�Sø�8pY�m(�x��8�/l�9}>r�W�PȐ@��
BnoŽ��.d'RHN<ox��>�i��I�G�5h9+ps4�P(�����.��7UUB�7�	(���Hx,��������`�ku%h'"��?���t��W��G�1�+�wEr̰TxiȤ�QG�+I瑣�K`=.��H��T}"&�x��x3&����0X[v�w������rـ5^̔E� ��$�R��[����Äqq�q�U@,�x2��ϭ�^��\�۞?tSJtv�Ack]����o�� �����@P{ۍդ圂he�s9"�M���f!�~�^��xD�~�=��?��t�v����`�-�<Y�C��������|T΢}���G��d�0���X6;�V�?������B!��=O�� ll<Q���%�0#]�×� fWY�]�&�`�)���pzY������9f��b"9b����!&a����e��?�j5����a��1~��?�'����p�3�l�t}�R��� 
L�D���ߵ��.8N4�ɹK��icF&�
(����u�D|�T��W79 �Q����O�>ȍ��+e[v;���y�ِ�qP����G����m9j�'�L��^�iC�O�Y��;�~c״��A-ڒ�Bq��y:��!Jp��px������n9��v�&�z1]�Oz�����|���0�*���;��U�2ʺ��ioY��0�k�O���x�z��%j#���Z-~c��`������/�;ro��#|�����rI�+wz,�ǢaW�{�2
t��� ¦��"�G%[@���QG��i�_N�e��v�z�	��A��Xc@	�>G�v�D���]k���d�޼:�$L[��5bF�_��/��ui���\�Vz�KK��L�⵮�8��﯅i�h�^YL4�_��͍G����$�`��ܫ�nǂ�)3��8�;"��f!���
|WEPP���iNmh���,&$�g�Jd=��i_�u()y�MSل}TG*>�9w��KѧF�L�L�k8P����Y��#ϟ��n�����Bs���*��i�I]��ގk��/+��e&�e�qECD��܄�]\�I��3��2(��w�� �/o��{Z�!�,w��4D�yC��-k�Q#�8�dύGዜ�F��p%c	Hr,a&�_�/
Eh�Pz-�$��bpy�) M�ۧ����źN����F���[�t��Z��7չ��Մ��g��\�q�z�k㾿�V���}��J����|nGIpK|��-�	���
�x������ 8U�0�r�)����0��kg+{j o$����e�(�C`h��KgD�1.�S�̛/���]�>J�^���Ho.��Š��|s�+�3��A�м[h�K�[tH���=���\�\����z�C�8��9��F����+;�]Nk�N�~lOoB6�ip⭮�_����p�I0�Ys�gzD�@ю�'��׍jBv5G!ۂp�^M�̴�Ղ<X�$����E\��@վ��Nl�C Mt2z	��z�SB��PJ��Jz-5��R������E�V.�4��&:�����#�!Yt�)�k3����H��ۺ��8�'�b,ھ���?
�h�x2u��`�2A�ʱ�@��'���q#�l!��zۏqVy���hZ���^��{1� �^�;X23�=EnyOۿ���0$��f@���W���7$�VMxE�~�ّ7��*��|�7 �j�B�d���?y�!��T�[���\5Qd�!�Sr�k%���=
������b�#��k|�4oM��/�j��6
��]��+�ak�|�c
ڵ��H��L�1k��h�Ф��\T̚&���s �����l�"�IOh�K�#�h0�
������}��]�)_�p��_��
����"�+{�ϙ%��UD�U;K�^���5-Ht5P֓3l����~71�p�bC�Ͽy�o\~p-�k�J��c��R�p���g�IN��R���?������~:Rΐ�A� ���on?��r,����e�r8Dv:��tN��p;N�l4%-��m�^�߫~&Dic�Ơ7R�KEi<LD���$]�3���{v�")���;�7���"cRS滙c7�2��U�VڿEGf���v9�o��[��l�_�e#�-)�ɸ��HLB��0 ��V�E����-d������hX6J�i�r�1�S�n)W��>�[l8��O�?=${�A?;hu��~�(|c��Ĥ��S���Tj+7��ߓ��;d"t,>���� �%��' P4k�~)~�2���6"�	�S�7�Q��Y�(a�/����O�r�Y���Y�y��c�'���EUx�L���!���	��o葃���l��D)��q�ؘ���������ݠ�����VIK���u�`�|G�˪@Rg"}
�^B� �P�)��|u��v^��ƥ�7����׋�ed���(y�5̶R���d����d� ���2�Ίa.jQ;��c���D�9��/��`]Ր��X��XTK;A��%��"`�o�(I.h+d�x!�Y7K��X���!J�U�\��h������y�#�a�����0�=��.�E��tȐl<���r�3��s�@T�4��3�2�M����� H|L�-��%6��8�q��ݓ�,���7G0�Y�i�I)�Ѫ�0���;��?�R��k��R�h��bș_�����׭0|}nS��S�dw�U!�|�n�����=�A��+ ��0n�]4�D'8�Ab 0?��X3��ۤ���Kj/��ܗ�(��[�R�t��i�Rm+ˏK.�11j��l���J�A��R��"o 7�G�>�+�r_=������JL�����Jwu9�al���puk ���;�!��y)�c|�+�+���{�Q'�3l�Da�j2,�C���W1~�.��RH/�y�N;��{��q "~�o�{ΰ2y
7�WȞ��	ᨹ%��Q�-"��b�x�[o�G����.rW<�H
Q�_Ln{UҜ p}�J�{k��BȐ�$�#�Ҿ�>jι��ţ��[�{�L���PP���d�L��Wz
�g��ҩ��b�>�V&�LM��k�t��=���.c_�{�Z���Q�"cwK�G\��u�0��
��0�hh!>�7E-̲z0���hXLn@������2_�^?��(��%��e���p��ʕc��yl<`E���ߖY^��p��C� u�����A=ݰ� �FJ�D˫=��~�f"ۈK���Bh��7ݬ�����8^�+�e�p�+	P.C�7a��+����R[>�?	�Ieq!�������҇}w��{��+�������D�ڽ����#�H,����"T:1]�����.~�<c��}g�D=�B|����������?Чe�N���&>��v�l��U>��HtN�s�\?=4j�0��dV+iJX�#EÞM�ί	&@��B��,s��L�w�G�^��O�54����`A.��ف�(����O�f�GmrAbI�ZfCn��
��p�Yh�e��p�Ď�)	�{JpZ��j�Mn+<��ܙ����>H���Ŏ�Z#|E���O*1�]�f�KGC���􄟦v ���:�C����Y�����3�y�����ؿ�^��Q���T��)�K�P��e���69�Fqn���-��Y\2�Ǌ�������g�����kz7<T���̉�f��q��^��$JpO��.5��h�{�s�h���'_��"GC�]�戭|�Vc�	Ua:��t�(�l<7�l1@�r��9��H�k>1w ����~�ͮFd����QY�c<����(C�*�U����8����D��ʞ}k�c��4���|��!��Y��A8�f#(�Z���D˄r ��,��u)R�ֱy�a>���iT�a���wq������`����4�����?`�}��{�V=��T�>�jeuSt)&���X4Ew�`oK}��.φ�=i�r� 9犲l ��q�H���z���Ƚ�M�o�@�[��`���Q�"��⛗f�%{Т�o��,������7�0s[yl��[+J���"H�U��,i�ˏr[�ou�h� �!���(�0'c�M`<�cF�v=���ߎ}ݵ����oH�ژ3�IOQs��S*�u�B��4��o��^yN��v�t��o#��=���,2m��w�������Dq*���=8 ��c�'QU���H�a�4:1�2�]8A(�\��d�F����C?aWUK�m
�� @QC݋���c�y̰�ÉV^��HA�_,E���� �5ށ|_��B �{��� 3���%"�L=~�,�o�<o�FJ@{#��*j�$u�ڡ��>�﹡r;ҋy�9�}b �94�,�*Q��[R/��`�Sή���9�}I y"%�=z��g*Y���,9,�U�l�x�c��#�>�}`���j~�K�'3�۟g��i�6���f��'E��ȹ���<nI��|��9����?���(æ�x��x�AWO;*��/�r��qI�D@Lq�{���[��8j����.���m�D���H:7�UH��
Xa��K�a9TQ��'۪-����F��yA\�]��ۿ��y[G�#�sF�(��w�k�iK����'C�y�#�=���'��lѵ��e�(4���ܔ�i$���<���?�	3�Z�k�O��LI<S�i�D<2��;�V�8�^�Ejn�b�!�¨�ƀc���\��&�X(.g�=�	�!�[E� l�s/}�#\c����+*[��^1��[���"r��zݣ�ˮx�O�/�Ͱw>k>�u�q��������"�-�v��O`86F?9���7�݅a2��k��6򘀓��[wu��z9떊��t����5"�H��\bz�4R�`Y8,lC:H��w�}~�Wʏ{�%�?�U\���_��Q��T�ĖGF_��o�B���O��6wV�i�ro��g��)�nجX��Q}=tk��e���Ȉ;f���W�m
��k}�hLP/�$�V���RWc��X33�Xi��=��ݼ,c:��m����X�Sva	�IQ^"Gu��'Q[ݻ�?6��C���`#9�ʭԭ_���	�7s	�y�I�e�|��'��m�
�e�.��ӱ}Sb��1Ts�d7����'t�t�/��d�gˬaj�vV��&����JFwx���j%�b��¿rcqv��C�~���a��D���G�A���iM��������b���l4�1�8%]W����Q����	�X���wa��d�<m��<Q}��	������&���1�"�:Z(�*d�`*���F��J���!�k��i/0� ����8��<0�ò]O88�VQfH|�u��z�נ�Q���Q��R�*49�"}��*��$��j_\���ad�)Lf��6e��)o���5��咝��D���A�e���5t�����vq���i���1T ɚS�s��0�������M�s�����֑�����?'�F��B,g��RF� �?�\*�E���)��x�;�-a��G�Lu�OZ\O���C8�b�Z�z&5���SS���j�)
��	q��,����]��V����)�<�΀2��RVCޅ�k�fR)��	ؠTg|#8����t��*q��;k9h8�8P���<�+Y-��k��+��/�����)�]���Z��B���ZO!ru����i�P~>�ĭ^���+EֆP���::]��զ�u� FJzY�L;�k36U�o��ֺ���x�ZY��;�0�D`�W����h@���g��� �KT�tb�A~i��?�y�ji@!��=ޙ'���+�Q�vc��&b8�wJ�ב��AX3^�2nރ�� >m��)I�4�� �njY��<���˸,�R�� ��$�vD�6_#�ᡟ��:t�WR6�|Y��X"�[�r��0��^�aa�0D,�/_�U� �e{b��GI��V� <[��2c���-j���5L
�@Q��{��=�U?*���)�߃����(;CJ7� ���懍{ـQ�%��>�y�kG.�Jo,���ByN��H�}C��ȼO;��n7M6/do[��&��.��k,cM_�o��/7���ڋ���#`��TV[��9B��6�^�N��U�>0����r��ʚ�ߡ5� �u"I�O���2���4��Sam0��6$�A7�JЂ�Vt\_~=���)����Y��\C8L"�^+���U�:gn����h�,��$���P�\K�G���ݴ-W�Y���9yy	���?�-��!	O�t$D�Z���^��U����(��Dk5�����_��t�4�x{14�(�k$\��c��={k�j9��ԭz�E-";D�UJ#��2�JK�F����7<��MbJ@�9���NP�F�;+R���J\mVD�l��Oja��)w?��`��n��#�,����T�(&2���s��$a!XLڐ����=/�xT8���Ok��}W�Y~�㻺�)�Z�E� �8�̱�\'^��(lc'e?L��3�y�Wb蘔�v�����%��վZI�8�ᇶ�)�����69�ٔQ�6y.s|���<hSۂ���̪�v�?��-���礴Z��hģMCχ����7���D�u;@�5�b�`	��~�y��8����q����\��m+�+hҰ BK,�c@�]�W�e��4��Ɂ��Մ;1?���w�A��XZ�k�͌��E����#��v�=�VU��C�w�̆\��^1��0 q���,�����f��\,ܽ|��Tu�V�X���z!�.�}'(-�?����H#��������A���ѣħ'}%J�U+X��^������C�m�(]�Th���vAs�"�-��
�H��F���4�"A	���EK�Q�M�_H�bM���D�� ЪY��Wyײ��ޣP[�����;mN���?��И#��	�l%к�,�p��θ!��ز�|U���x�aZ�([�1~LI�$,ycT�c�N5�7��#�N�Z64�k���lYL��F�`�	](���	�~<F_���L��-�����#A7��O��D����/��B�_#��pZ����C�W�
^�h=h�^��3�� �c�Ä �Lz�sþf��a�����Ht���7=ǁ;��b��8Y��N�B��8)!Ѡ�F4}b{\�*��[Rj{�� C�&#�����j�~8��h����z�&=ߜ���b�N}����/�{�w���ݓ�p���<����P6����c�u�qP�сz���V�Pm=�5� ��Sgn�DFC����ѩ/���D��̌'\�@��'�m�T8��Z�:�<f�9����o�3�ԏ��~��r��é�)|��|MǋD	���<��9Ad�ܜ���[�S�#f�@�5�l���.�< �ҩ_��u��^��u+se��Y����x��50�������~�z�����8G�
��/-+�۷�}uw}�H �l����/�����
4��l@~���l&��� �RjlM�b�B�_��4B���w�i#]�iH��Bij�e��U��@Ϥ��d^-�CN��9�h��H^ZA) ��r�5�dzJ��",����k벀UA�7Grq [i�y��%�^�¡��5���eO�W��G�)xF.A�CD��Rm�%(�}n	T�p /¸/�x���Q�t�xɄ8���T����M���f�����l}�>����]�����fCk����fT��z��z2# ��M�^�Gq�>�1�ru���r�}�&�´6S[�_���l�!��?V�p��2���Lm�z�@&jg�f<Vd�T��M>ӛ�T��t����!�qi�����U'��Ћ#�gO/K �W�ynXH��i)���U�9$��62Cٗ�\�2a>ڈ*�Uck�0�I�e��k���=�K�~k9^��p@F�I5O���STB�MN�jOC�G���� �?�`W'(~�����������ۛUU2r)��3�Ә�\X
, ����m�n�ad���q��f�-��3E��˩y�oSq"[iT_���4��k����������o��iD�1�y���n�T�Y��C}b�()e����6>�\�I4�!��Wn��)�od?��c�����"��-�Bl�����n�����b�*����Qu�m5���$�>{p�� �jվ�=52�J�r�߳IWT*g\q*�2D���B��)`FI2��T��)~agLH����������h)�ԗ����xKS�O0u'�������8�q,o�A(v^��Pv�^�0/_�Lc����������<R��c%C+4_����'�!��B�v�*l͘��R-F�<ȇ;�~��:�l��TwEJEؓ��,c�N�~�+�e�7s��~�P~?�f�yG�Pw���ޞ|�!�;�G��_�.1׮-U��'���~�(���G0��n�8�����UY�W	����V��P����\؇�bŘ�0�`c@y��$r%��S7����gՎ��}8�y���-hh��5~�s���|!���[��c�����A�W	���@&S!��.����.�x{@��U���t21VŲTP��� 0YO�7�����詀�,~��:�D���=��{�
t͌qA�R�k׆�d\]p�%��t����5�=��ڴZ�2��9���G��(�� s��RFt���A0�/�EV�e�4G)��4ˁ��)5i����a����qf��(��[��"�|��usUgb�O��hY���������a�յr�t�$�E��:�"WS��:z;~�G��rz=�~u�o��xsH4ɷ�J)Ň8�3D��s˥zsi�r�Qe�(���`���8oD<� ��ف���J�e$PpY���V��pf(��<R�h��������+�4@��bvT&z~�˒���;j&[W�Z�lC��&�nop�|�f,�J���ȴG��9n�K�/��ˡΒV9����v� ����3GAR�8��ᙓ�O�Ȗ1�yL.	���j�"z��_��z�+s��cć�Zh'��C�Jyi�H�DT��# _�\�_{T(=s���8DR��P7�P�v���V?�odf��.��T'?���.��9+����d��$X��I����H_��:.�	A}
v�c�9���`�,tJ�Ðy�E�.��Y�<���AR	�$��d��+�ܭ#��M�b���s���tr�R��\K
�[�>M���xe���Mpp���NJ�X�N�=P�&d�'&U���wCekܱ�}�G��;p���͏Gu������w��L^���;����!k-U�`�|�����E���9M�����ϔ���_Y�i��d�B�L�1_���Ov{��G�5�,x��Y�㫢J,)V����ùVY��a��HL�ˉ�=�,�$[H�G`��4HM�r�Sp�apF��A�'jYt=�c���S�^�#���$Ev���.�z�&P�i�9�����Ox�;p'����L�W�L�ڡ4.��Tl{�A���m�.�|N1������+���
f5Ϻ2��}L��4�ֶI0�5܌��9J�a�U	�~��Di.WFU����q�+�#�Lo�h����IW�t���A�!�b|@�����$$����k���2`#�V��&r�ܳ�lߞ\<��H}�e�=�N��c�����҉�_�0:�T�)1���.ȒD��g����ޏ��"�n��E�[l^f+��DY|MG돡2ZMWXt�#�·ɱ�=�e�(��BL�0�� K����}��C1 z�Zn*'i�50�#)�P�+�f@�P�z�n�'_� ��4�1�D#=�(C�������*y�.���8�Ӕ����� ����;AH���������D64��G~����z��p�����"�w;꫌^��{*��EK��BBR���W��t���h<�Oq
x2ȷ#�����Yx��}3��x�����2���3ht����1E��Gm5�9z�h�� &�k��M�J-�._�'��l�^��=����nK�Ϊ�F'`M7jwFr��8�T{6�������k�׾+�T/(D���vm�6{E�G�
�+v�L�R�X�d<]�����J0�_]����j���1�����l�J Lр�AO��$�v=�>��q��r��#0�<�~G�y�&���M?TAg!�,�[�C��On�AC�@)�Z�&τW�_�V�T���ݿ�O�A��\l?�[!]�ޢ�2S�UА��0e>9F�9��d�c(�nl;y[2'm��3����k4���L��	�����@Wj���$������j�Y\�S�x�󸬕��1��N(\���
F 7!iXy*���������`����������g�oE���R�CL�0<`L�Z�pw����Y*���̓um�4����h�������3+��5;-	�K�VG�� մKc�7��m����>,q���a��3�wc4[a�(�߯\�yH��fߍ��WI�W��5�Q�%��]�:>3`'����m����S'tTy�̲nv
�z$	Ӂ`���T|�vɑ���1�y�rY�,vV~��'p�Y����}dS�φ�.
6��	�'�x��׋/DR �L���8�侠��L�`E��DyA=ƛz�ئ��c���~g��(ň��p��j�XP��~0}������a#�`9;���q+YK/ z�h�`�~{/��N�n\������_K����ԓ�D�rN��G�����N�kOe�<���1kD�������4� (����{��7cJ�{}Y���t��m�S-��DW�ZZv� �:.-�:l�G�����r���s��f<��xq#��Ϥ&@���%H߽B�MK|?2����u��N��j��T<.2C� o	.�.I8���f��ZJnO<��N4B��P��,,��<�7������zs�&^H��r@�ͻ�����≕ˡM9^�^?B�X� ����:h�t�n�޴|esM5r����:;�0G{������:�F�������Luot0~֢V�tP�@JJ����*:
�bj�	��U.�`\��ߣ�$W{��C�pZ$)��ß���\�$�,���<�ݞq����ƨ~dR�K���U:�����}��7o�D3}�v��;�u�^�򘉧��\E�"d?Ɲ3����ϡ�J�.';�5K���J%##2ݏ������wC}bB��E�*�'�z��(Z9uS�noH��g�T�6b�k]�����G8W�
��Iq�F0�!0�D6��;�����K�K��p�N�T1����0���2��a�
��X?���L`� �ʜ6�v$���U7c~�Rou����'eK﹕������6��2��F/blʻ%��(��/�%�H�k;J�,u�Q�����#�D����K�l�
���T
R�i��KB����U�&�/�%�,X_)��مL�G�=�]���N�
�|R#v���������t�� �WbkȊ3C*Y��f�XJ%D�Jp�L���A�?ԑB�{)�yM\N�`}/E����B�L�b��^3���x�&�XDR�ߪ�/InC���	�k�n��c
��Pd�"���M�Fu٠�>�X��,)��d4
韎U��J�Eļӡ�S�`[��[�~S?����ҴlV4�D뇾�.KT9��2p �q�~[��U@�=֚F��M��,�oV�k�}���jA�q\��=^�3�R�N�W���$���]#ĕ?��B��~��bG�}p�L��(ϋ�t�I��έT�y$$��h.I=�ӵ/�[�
���(3H���\S֪@H�M���?GX��((�n6^��X�������v����1��L��g(dF��_*���v)�$'�Y:{�p��^�����tj�ĮN�9C�w�k�L)Q�l�4o��z̾�^|競��rd~��ƽ(DC��±����2�"C�S��4�~WH����J�;
��/�մq�a���.�X�ē'	�:Nf�!!"��K
>�	������XTɐ+���7=�>�'����we`�� ���>BA+D���UGɋ���V�u�P+��%0���ѼR�7�X�u0���SK�C�c|T�B�5ۚ�ye���ڎ/�mxX�YЁ�XVaA������5R�fr���	�i��ʸ�}I��ƺ���bh�����E��&M~j^LEЖ7�v���G�1�k��j���d{��{���Rބ�`��a0��;�/M��~P	�Y�����K[�>)���U'ʡ��n���㇐�>��m��k[��H�_��4�+�<�. EQ�5�#ֽ��6S�3����oD��������LDA�ʪѵ.60x�``�l�l�s�y�҄�a���y��2�d�������#}��,�c�I��^=!�w�����| iČ�?�i�k(`Z��%�� 	�(D���J{lk��u�?'�-,_�)���"T]7Q)i�ap'+���vE~J�rA9�AU
��s���ջ��2�O܋W	�-�N"	�s<1��R��W��~��^K�0��P�k�q¡�L��Ρ��9'���}�����L����^@�^�7�n��hzɗ�~��;���p�"%Zk��$�:�Q�Ph��X[�|���
#��wBf�3or=�?�X�X�eFxZ�/�4p?�:���h��B�Ѐ��*a�'H�gBo��D��:�$�Ӯ A2��gm���ɠ�TT��<bQ��4���k�,��os�S��n���j Xc^V�K�����,���U�G��WY#l�\�}S�\��1��b�<zt�ȅ��зLk��cL��59'�-.ڽ� ??0Uk�����bdd8�ZS��]	��� ��k�%,_ �zp�1��G��5,�D��N��[��v�J���=��9��,�U�� ��~6�c^��	�r���������4*M3l��$:Ks�4�9DOKb�D�=�wQ!Ɖ��L���c4Κ�Rq����mE�]�U/"��ɝT�\�K�RϹ��%+uKǭ��{س�T|cI4���~�W������z���Ujw��+]<Yf���*<p�r��a<�����0� �x��Б��N�%1_H��nG�r�c�E־Y�K5�x�zhK-���T����w�����13� K�����wً6e+u�o#$�������JMn:s࢕�2�s��������@�;+T�T�but��0
�=��E�R��/r�u��:)�~;���r���k�{iX<j���*-�,Q�]|n��""�G._*O��f�����ˍ*^'J��Rh���q5h*�+�#��~�M|I��B!��)�>�H76�)�R��'���� ZC�axw4z�9�~�3��M�����ី1ru���HYwS�k���[���lEX�4וְ����&�#ٖNo����s[�v#`95�Y�3l4����n��5G�.Mk�����ɡ#t֤��=h�t�ڍ��a����A߁�RJg_�%�_{�f���_��]��|��c4�#��s^漜��U�5D�r��O�f��"@ّ���Y�Iz�m��U�P�,� wp��)_��t�aa.h�lKdz?}��HP�G�H���I.ơ�����1,pK�*b} �P�l��@�('#7��� vW�J &��q~բ<��h��B���L���MFgz]��ә�0 �Ė9J�l@�g*��9~��Q4����8D�"}��7���w��&�I�!m7��	�;���x�m�@c���r�.����6Ìo�ڒ^쐁��G����'�W2oEV	";3�n7W<;Ӎ5�lx��0�h�����çp�5x�}�hfSm���'���,Ȳ�4TAƩ�������)ߕ}|@�y���
͠|�'O�R�'ş)jnl��y2LWe�҉�O������r'�H�L)4O$�;�:88�N�4v�q��Ù��@���ʐ�GvD��kЕ�Y�oi)�\�%�F!����X¾�k*GsQ �FLF����o��E����2�BA\bN��D��[>��" �} ˘&��=�jy�W&\�OG2'H<˦�8��s�Gv����ط��} /�r#���)
HgE(i�%)�t��ض���nƲWR�ț�t�5�^-�AIWQ�⓺Z�,�^����/���2��Ts�j���R?��� �8���&΄�47i� � ���,a��a�`n��ڎm��~I�mi�������I�g����k���f�8P�~�N�$��h�l�t�B*u�U ���W�=-
�sz`3?X��6�����C�Ij��n�p>Æ9 �sm�R�,'�%�B�j]��kz�����<��.�AFZ��L�@�:Z4�~���F2������ē�j�j>`�C� �-l��V��I�1.�=� �t$��>�^:(���N�:�U��y]E���96�����Y��s����M��߱r�\ND1����KL�̩�7�H����is��RefO����	����!��K����h�3&dh��s���E�F� ���R��C�b��rڷ�b|��K��TZ,�@���A���G`Ƴ2;�������~�\(��Q�l�({��EM�w?8������	E� 2d	G�>�~C���"F!�M�6t��F��>Ms�ɸ�D(�����n+5����U���?e����ܰ@���*MU�d}�+a���:�лP[���F���O����:jog��<[�:I�Ft��]I<V�<�i/^�mxǛ�`�2R��z�� D�^͗U�G����W��6�kbPv_s�2>�BBD�C3���g��� ��� ��7:�B�}c���$���1�"�9m���Pm��P���G��:?��)��X
���N��{��ԋ8@ΙVv���O&���Kc��h<���0]�[.��lJˇ0* >]]w�!�RB�X��8M�3�+� �Q��'����^<W�̘�򇴲�G�yx1��1O�F�>,L^a�Q��w!����45�G�s2y�����J������7��%��əφ��c�U�Qy,��96�5��
�շ�Q�����E���g��D��W�%b��K���~�G�Z_Hʲ��G��Y�mY~46���ɞB|� ��<Y*T�F����4�,6Wn�=+J��4c��7pB�m�3.��a�`��dЇy+<���/�L�8��ngTVr���@pd�؄�EW�
�A7�@q��J.����z4�����5P���
�n�M�/�#����]�5�6%b�ㆄC�K뙉��c�4��e(��NP#!�l��<-����bJ�	f��S�{������._�bFp+�WX��F$��bA�i��N�V����5��)���k�ی
Hp��8�V���G��t���q��Y�c�-J�HH�xu2�]�h�p�F�A�
�l�J�Jʫ�|2�}�SCHkƴ4<�Y�pM�{|��A1,�� j�X�^���*jT��:q���+�MSW����0�B�TYs�a<�7�=?����l�Wv(~��U}� ������}S�M4�ng�+="���X ���M���Ц\�'q�޽�\��It�C3Ҭ�R��9>I��Gp��=5��"�ٸ�Oaj
�P�8.� ��K�K��lקHh�h>��5Uڇ3�{�M�;�Fm�P��
V<�V�$�3�?�{�����;�_gB���߈/�'~eW(� װ�}�p�1I�{�Jn4�*����۟���w�A���W<�gT}�lT�!E*:�U���ݍ�����J�8���=�c�[�+l�o3���|�u.ӫҨi�8	�y���U��ыS��)�	=��ьl9��o�ƹ�Ad$�ru�/Vx� �ms��m��t����Ak|-�N�2�f���L�oߢ�N��{�AX�?2�5
���/�����X�-��	�$I{$�o�z�Y�R��hm��j��s��Z�vB���l�%w�꫸���u����D˵�8�0�ߚ��0V��$  pS7��!t -/��v�\R��~����6ޞf1V��y1̱֒������
g/���-���� �iZ{��Q8�ryۧ���.��%5�"j_�J���'���x� ��{<��@Z����UU�Ds����>��CE�5#;y���^�#S��Iˏ�]��9@°��ӳ�7�thzܒ:ޛ$@����Г|��  �mx�{���"���~@��%�[-����u����)z��O�M^�=_?!�jU2�Y ���)D�B��vJ �>�<��Q��u�}��ZV�՛��OJ�ۯ?�UA�3�,���[ J=��S#��hb!Ax|���;O�Ő=|V=�.L���yk_I8[p�#����{������S�1��ERr��}�Z>����Fn3� ;�R��;��+�9��末gΑq���}�,�ΐT���/���T���� ��f5f�z�d�Y%�9����}�(�*AZ0��*��؃�S9��c`�fh����|����؋�ү6wq�.X@���<���P
�pCm�K�����/��f���\S���I���a�tλ*Z�;�5U^��V��X/9sB�&;-���Ayy��l(6s`�]�ҋ�AQ��)K� 4�>T���\��1t�C	'g��p�}�^P�,�)WJ4�W�6�J\̵u�����(g�l\Ө;&����6r�x�G�p'��i�ߥY.o��?nde>�?�"���� �k����!�l�Ó��Q�˗^��n��RS�3$E8��m���yU`8>\	���Oqn�Y7lΘ��8h���F�*sCl�: +��
1�#�q~�l ��q�;���S�I%{pa�d�3�� �N��R���L�|����75��HP��#*���G~�3E���a�<�3t��T:��?�y_@�����Z��6�m_O��#�}`��KlH�F�S^~{ze���hX���%r��"#�=�]���4�����e~T�ۼ�T��q"���$�P��e�zww���˦�pO�r�v��j:"�F�}4�Y#	�ƴ=�!�W��}�����i��e0m��p�Ζ�J�5���r�C����t�EL2�ίs���tnS�I�+��)>,'�G
�E� ��NJ�UziJ�����(e��/w��BN�Z�������t��ph��W�ޛ]�����ˇ�	��Ѥ���W��tV���s��H�5	�@`hq�+넽F2���-��Mb�AO��Mُ-��R�oߘw
�w��+&�� �y�b�%d�i"ߜoSVހn �DT�xp(D�W�T�g��U.J����M7���Mk�<��o�ޓ%��׬��"�%�1
/H���e���g�we�ņ�ŏ� [���)#�8s}�-8 ��\JL��ƈ��W'��ȓv^w���K�å!������x:�q���#߀�<�]R�B?�P�g��U��
��$�\M\���nOm�J
6V�n0H���=3��R�P�&��@+Jk���(�|��tZ$���\yp�g�A���(��Zx`�שF�g�ɫ�Zq�l�lU=�����ѐ��MY���L�z''�X���y��+���S�ы�W��U�d�oP�Ѫ��`v�Q�7���d�����!��>9�<������G
t�!��L���@�B����W��#�����+5�37�)���p1Ƚ���=�~~�a�f�9�T��gA˴ �*�!��F[�S>�Q�'��*�U��JJ�����"��Β��z�����8jޅ���O����U�`T�g�uYt��5�b�%���}�:��o�9�j}�>���{��CH5��I\�����#��\]Z�CMm���;~�����$�Dݮˣܷ���L�͋�E���P�s�olyJ�Z�]�-�U�>��#�C�dy���۝�q�K�z`(��PO[ ҫ�O����V��-�[�|���$��D�1����1N4%��Ot�V� j'�?���)��,����B3)��.]3�*��p)��n��#9��V���CNgN)��]b��Z%�ވ1&SJ06
{nJ\���/V�OW�f�P�"X KɁ�>����B��ۋJ���'������>"^�#���]���_�3�?��U�Q�6�AR�䘚��_5�O��5j�]#�#D�c������-��</S�d��v{�:�Q���Cj�,�hĉ~_�rx,�;�!��M�ڙ�����(�.6�qs$�˔��������5�U筘�Mx������f�p��)`��v�3w�����tп�ྻ�&��Q�=F9�)����bz���WW)[0�v�r(S|�n�zQ�S�O�j�e��(�(Dɓwu����-S�K����>J.��_�z(&�
��|�z��!��3�a�͏��\=UX.�}}39ʝ�q�?Ao��T�0�F�1~5���T��l�'O�f�[UAC�xߺX�z��/�ңĀ�]Myq�)� ��.��~�&" �B�n��a�Y�6��
���:�Ҩ����gU� %������K���2ʮ������5m�!�K�w�����U�#Z���o��'�4�t
��'��-\_b����Z�z����d-a���g,7*���*��縃����D�M�C�;}+�-S��δ����;�r@T��!�(��"W�٥�����z��({����$5�Y��rB�2��.�K�.�R�[i�{�S��pٸI
��������+�Is��V��->�4�¡�$&�-�� �T��A��gc��1)r֞'	��	�uR�J����As��2��	)]�Z��v'r�Y�CY~�ԝ���q��c���P9�{]��sS�B��.�S����Y��R�V)se�`DiX���
2������}{mzAi�g�W��C�mm}�Ѩ�4
��j5ӧ�:[V��$�r���SJ��މ�kho�?Q� ����Ae#�R���_�_v�ك|�3�m�w����4h~#t^V��ך��R����@Pф�I]�1��Aꩿ�J>(\45��/��F�-��4,Nŋ��Ӿk� G�s���=oѯ�F��e�YZ��߱<����,�����C-7��E��K\z|�:�Y�����u�C*�90�ϟC��g��\�%�s�+�>��F`�a��X&#��o����E�H#�g�*=[��;Rr��"�Z�h�Jg?p�`�(��_��X��X�W_�d�ݍ�� 8�J��T�v��3�	����N~E���݌���#�]	� �=��(�z�}���Y �9-b�)>Y��ӻd�p���;�a�	�L&\�l��W~�hbYj{O�Y�=�t�ťS��L8@[��X��OwSsW}�:�ti�(�d�o��m��P�#KC_�J
�<�*h�̒0$�LX�`���\���4��H9�)*!��������ӣݴ_.�봟�9/U��SZX��_ӡ�s뱼+Wf3��Z�s@�@?tp�����}=��tk��H�&h��ۦ��$5[c߁��(�]�.��7���&�v��"`��+�茧�����R�fD�mфb��.U��f;��*���89�?Np�``���+��Ze�B������"�M=	7�'�Jf����kDzR�`��!-��(`ӨL~U{��]TC&X[��C�Z�ڙ���W�����`�%d{���eӬ���"�8Cs�]��51�2�!h���I�#�vNR����%�r�G_�Ϣ�O��L��Mm1!8���ԍ����G�b���z�R�^[ՋP�	�F{����
k��$��fXU���qS�:��K�ۤ�#�_ؔ��Tz` L�ϩ(�%PL�O�m�"���v���#�#~ N*�tI�1�s�M2�������={�S�ݠ�pi�ф�P8�.%���]�c�;��2,�F��`�,G�#�5���/�>�I}$.sY��i�YSl�����BUs�����C�`g�� �������a��l|u98�O����U�s��:>��`�뛠$(>I�/{,V���n�������΀�_�v��j�
]�V6F��\��A'~����"�)��+�!6�4����1S0�]�Ͷ���S��n.�6�XU�%3p4��w�������h\kL���*n8�`�!���qWI������J�m���ky�3���/a����!(����p�[�C�5�άQ�G%F�����B�.����VC��P�rI�s��1�:��i�B��*�u*����^J묕�¥�7�w�$1�R�p����"/7M�s��م+L+���e/ǔ�[%n����$[Kqq5I&1��Q�(a��ϻ.�@�(m�}-=I����* K�X���a�,�G`�>��NG���Ys4.>h�M���ф���Tϝ���+���X����2Z�=^��Xr�l�j�&��17�)(�<�jgvU@{!G�����a��^�`wo1����*�"��!]������/��S}�������*�M1�3����G+U�	L��Gi�m����(i��v�"�YQ!�E���T��?�}�b7SqJo,{2ͧ7R^G�v
.=��_�,V{��b�ۣ����O��1ʗ��|s�@�<�u�z�q� �ȳA�T�N ���v}r����qVRl�i0ԭ#�:�,~�NVi;k�s}גQ��)��jB��l&�O�@��t�2��j�ʅ7���$Y
��~��K�Lt�^�+�m�5C_y����ܭ�k"�yN�/0�J	�O">D(0�*�h�a� س)�%0h��?�a)#�H��+4_k�M�p$@?88��Pۙ�O`�~�s���v������u�;m�%�Ft��)�Sp|��t��=R�l��äÃ��HJ��`�����'�Hl�dڡN?�	��M(�Dݴ�A\�}��;�V]�[1�$}�S���d��x�����%���3_��
X�	Z��m{O����'�R�K���L�1�8���J�8#����Nt���u�<}�tD8�F/���K�Tu&%`z33�B��]�e��׿�.�"��"��tS�l��ry��_��hJ==^�,G1�ֽ�90�ze�8>� p�^�� �i�/�c7���ѣ�AG��ͺ�'$����iңm����D��zlgy��L�S&-������J����0:��('��f@L%�h&����� �6�W�o������]㔇�ʹ�����}�����?)R�	���ؕ�ՐV��<�����	��q/�ᩁ� 𔜍��1�D��~��'<�� #�;}:_��H�{�͛NBC����R���#:m� �!������l,� <S��ٶ�j3KFX��:���|JB�=*��""��$&��z�{�$�Jޫ�>,���*r$\VD\0/���>�=&��ߺ��(f]�^�`��C��u��I�,�Fւ�?M�vCLEf�I.}����]���\�#�B0���R�z�"���G��9�u܌ ��W̶������r#*B�/��kx�;]<,��*��K�r�P���T<MoykH��sQ�6�
=�ַ�F��$� A�Vع"���}�|�_�i��a���z�W�0�(�Qz�7!���k���d�IC����C��~��ͷ�m�38~!z��������*j4�ȣˍ�ݙΐY��=.Wf!%0p~kά8�^����/A�8�Pݰ��z��k����wv.������q|�"୯��m���02�K��'�����BƩ�Y6�/[���<��o�H��H���@�]
0�poF����;��>(mh�7�I�m���+�����dz������Xjnly�MxR��iNn��R���?�	m��;�;˕6�������������S3�K{���B ۾���iɪ��-;A :�T�	�+�\���y�R��1��˰V�KՓ��U<��$�����QAm=]S���q-�,&@��n�BH��g��1�-?�J=`؜F�拥��^�K<�r�\ښ�Fyz�%?�j0I�
�����2/Mk���s��x�&���6%u(/4>ի�Y�1�������!)�3�7D@ɀ����ň�V��^E|�� ��̶��t��W�6� �^n��A�!b����?]&�s]qin[z��8��6C#>�;w	����%��<�)�FLK�$���AX2(�1k�r_<��[�#n%-����I�A��G��k��b�����=^)t�v
]�n�\������f�K�,}��}�"�=�t �6��a�b��?ǣ�f�Z5���D���A��
��[9�ntۼ]���%+*���T}^йt>PU��R�X�,��k���m4��1��4��`<w7nqP=ʬ�� Y&'hN+� L��f�4*c����70� [;(��:G����UL����}��mkp����`�y�j��S�C�6q/���l������r�k!�x�~�׀��qz��E��I��������s�ҸDKq���[�6�����O�j4'�1x������d��q��U�����kA0�
���KM�Ex�z�'������n�'=��y��A���1���+.>=e&���!�y��B,@�<��q�-��()��0	��'�:ë���q�|6"M���$2c�a
�3ny1H3����Yr�IΩX�� ���
�l<�O�%T�Qj���ɠ��	@���{:J�m�F��� ��h�]'�����ؗ�vBA��g�"�>�����-�/Z����m��R��-�B|J��R�jXRݬ��ČlYĪ��I�P����������OT�Y$�GVO��|H���W��њ{�%�"�'�VwFI��4�V	h)
l-~m	���"/vL�pj
�h8b��ޤ��b	7�W����2#월��0��l�s!�n�T��7�	Pf&6��@��������z$�ѶU�;	jM�u}���hy�������/�q�z��%>E��fڼ}�&�7+J��b�Ѱ;��s-O<`>��������جv}�W���%W	�]'l(��,��q��dA�A۴� "Mc��e��NmO���'�Vx��ɥ4A%ɔ��K�f��}��y�4�4i�E]�X���Ɛ%DL�}}X�IJ���PZ��o����߳o��!.Kn�c;"+^򩆣x�.&�=�Va8�{IM]'�4��w��&쓿�R|�����PWF~Bqq�V��i�5�X�Q��hH0�T���B�3��Y�Z��Vs���@i���"c�۳q?��R��Ӿ
�t��� ��Ff1��uG	�,&r��zaH�,H�Z�WDظ�:>�*��[���U_x,]ԓ���~���Bl^,�%9�pZ�k���s�I[Z�Hg��0V�Ms�O,�oX+N&F\�H�q@��G�V�J�Ŕ�ױ� ��DC9Ias��/�n�I����KP�[�����3�)9&?ddt�J�`��Y�����x��eg����v �".S�Th�n��7 ��g.&�(=�� K �N��\W]�%65B�L�coD�|*�
("L������!���憂�[qx_�P=�4I`���\���P	ѳә+|�ux� ���k��/���xd�Bt8�2�P�j�5`�
���Τ��'s*q�J����9(T䰋8��������+f>7'���U�i<
�|��W��pQe�6�\����as�4eb��5�*I2�j�Q��r�=uP�6�������3�qc}������Ùª�㾸��@Q��Y����"o^�����f5F*Ҽ�My�wspՁG۶vM�&O�����X�k^��y7�ϛ�@h#S]�8$�&qQ?̕��P�f����&��_L�x�f�т���E�*�N�0B��ƞR
9���=�{�s�(��>r8ӠT�������4�e�Q	&͍ژ�����4�Z�g��g�i<5��� v�W��bޕ|�U�kQsvr��Q�S�������c9ܐ�U�&�PBjOQ��
ƹ�a<s����!��w���"A����Ƃӹ����5�Y���)I�8	v�O��;�M����h��2�:��#j"K������Ԓ�G	/���� ���t0�ӣ'��?��z��ߊ�7ݴ��Ff�g�%�m h���dzu*�RV���)��:��Y���HyM��mfA�=���ɍ\�+��;c���'>�rfe����_��Vr�1������W1D�����O����R�`j������S1U/t|T~1����A�+�}�'Ê.j|����g�Z���52�P��S͡ˊ�)4�oߟ��i�d��;�"����}<��B��[��E�{5z�MK�`z-߮s�BKG"dK.%�G?�����m�0�lLPviA���pE���LW_���f�W�k��G45����3�(��(\C��S��`��7�e��Eۼ�Z��\�@{3�jR�.�D�k��V����� ��qW8K��~�S��^Ф��2p]��a/�{�d|�`�.iJ�5ͺ�N��EW��%3/�ka��X��FsI�T�C�W��W�I�y�
�\�|+��ys�\�5Xq�O;%�� .9_U�$Ͽ��	�m�7>�}>
�U1����h�����"�{��SZw捓S�C�
���ǥ2��5��0���(�'�D	�V�C�S��)���Ӵ.�GS9[�a]"�B�ܝ ��I��g�\�r�!�\��p��X����82����]��$�I;���F��b��$'���p�H�Ɂ��Y�	+|�È�ശ�T����!B?yy��VD
�o�������;�S-f���P�r0:��;�Y9�ځ����oc�����-��C� �:�ƀ@Y�=]2z���+�ը��l5wzc����(�ʹ�����I@�M��9�X'}ެ�t�5VMR�F[F���э�I\�	%!�@�V�V�N���	9/�e\�U�H�Hl�.��z�l� �Ib�)�|I7�H	0�����a)�[28����OB�=���+pٲ�X���F�B��m����M{�����<+�+����
��k�L�A3~�i����@~��;���p]�jvRi��*B�O���-�w�)'��4N��9Id�Ϧ��0|����V<���IZ��b�WD�Oz���Uf6x�ke��sV�I�P-�f�A'��\�P0;N,`T�ӕ^��U(OF�!o��C�M5:�{���dZEaaɑ���#���E��&S"�����?�r��w��Eˊ<]3�#��A����1��Lx��`���Ҭ�54�!�d�f�p�K�b�)S7���WܒrH�g��k?�\aB�H�fx���s�Bz�ͻ^@�7����[�N��)�h�-�����T�z�ݬW�4� �6t�$�)<��"?�v �v�]6��$�C�i קo��Ľ@�oSQV�7�*Kr;l����f�+�yI���6����^�e��0�`�FUY�o���`(�׳�N�\VU:�E��a�f���A�=<��G���p&����,r���[���=���bG��\��ph�k)ڍg'Lٰ��㲱�7찆�A]]XЎ���bO5!ꔤ2cZ]�v�T��f�{��a�M:�?(s�9>,�I��<�Z�<#�L��\�ld �Jv��P8Z�!�84t��7)V�`��8r=�rR�W�l�	s�Vƥ��3ѳ^��)��޷k�C�& ������avtZg*�~����b���T��>����N�x���:s���ZJ"�2���?'2l���f���+���~�h��c֋)�>��/�$��],2{�<y �-j����ȏsΆ��.iN���_����>���s�v냋�� 3��I*��欕���8������)؆옕5<��Xc���#e�K��D�2a�I��JCi�8ɯ��E6��{g��Џn�:L��p�E��3렻s�@#���7�HCve���#S���F���Q����ӳ�Q�&����^����u�;��Q����B���]4ј�W?�>&b�AJ)���a5 Ly`l�S��ߩ���I��7&b)-45�����kU�3�]0b7���uT,/�1�l�t4�a�`�#��\��]�� �m��� ��������F�W#��I�L���JN$]�ͽa�1�9b.��f��8�.�Ҽ��B����T����~v�]�M����6f9� `��-�1�j�5�M����I�(VM]��^������k)��P�.¢"G�|����g2c�� |{L��;IAĿe�Z���2�Ph���tħ}�Ln�{9<�8&S�)���1�KA�&a�7�B������ʿ�K�Oh,�;6*�/��պ��tl���<%�����+������XU0a�?���[s����ȥR@�[�:Y�	��}�F