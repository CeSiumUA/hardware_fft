��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��������n�sv4��%-gϨ��hd_�K��f̕�9^T@-h����i��%F�V���Q�%X�q��;�Q��l/��M������Z���ȶ<(a��ك��BXƩ���<�L�q�׼�|3�Ee�w�/*�������pY�V}�hiF¨��}��ro�Iv�A�3zc�ܑwN�8�g���sE>D��*:J���o��Z?������R�:Y�9���Lޫ(�{;{���4����G�Bm�G
o91�5Kc�����'��+��˞AR���w���_�҉��T�
is /J�v�~+cԷ�3*��:�c54Bto�/{v�1oh�:���np�x�������g�E��գ5���~�jO�+�yX��+�2��APn`�}�q :������z"%��R�v�ۆ��v���i�'yU!�$q ��ٺ�$z	&��m�0�QomVP\%ڻrC#���k��K�bt�9か	�}{>����ݑ�s�<���>�O�K���޻~H��%��Mq��N���>�Meo���\ت�5b�U�g<#���:	�a˕/.rJ���1�?*�i�n.�����W��7$���t�x�~��Rj����3� r�Q5�tR�#Y�A��ڻh�z	\�A��ێ�@���7"�D��A�U6y{��"�(cUTB�.ϫ\]�mF�d���~`
_0Ɵ���<���Z#�)������$s��A�pQp�l�%B��P��2��mܗKnjYAA��y6�
�iCߏ��RVS)u�veD��k��Eƣm��ٽ]'d=ހFw$=/�w�׮"�E_$�T�+�M=�R����~Hd���V��8�_�LZ��"� ���h����?263Z�BI�h-lֵ��@0.�e6w&vk/̏	�j[r?t�0:�NAU��r=�ڈAI,�|�Y��ȲP��K�0i�!�� �4u�?Fx
�c����j�<W�dȴ�ōqc ��;�x��m�i+c���M�=�p7m�φ�1�5�_��+����4y̘��' Y�Ä����)P�N�W�o�]������Ա�D�r�	5�G%qC��='���d�� w��PRÍ�%$�qP�׈8D|���ݴaW�Qi	.�zj�s��i���wo��#�f�q {!�B��DiA�6���VB���YD ��oZ�����:��/`0�Ɣ�;�5I���6Qr����ԛ��q���ڐa�Q�Z���1F�ݰ������~O,��G �a2�YѴY���K��5���p�W�� ����$��zA�ĸ�:�����D�{R%3��Qa<!��
*v���8�#�b���%�C\M����	ع�[	��a���v*5�p��)T�� C��kܥ"z�uN����V5��J�~.�� �U�v
K|ӱ�����/�:)��E���6l|y<td�������&�dّ�����ϓ�T�8+�O��X��1�Ґ`��A�{" ���/�Lf)q��eE�Ӻ^��$����$<� ii� �,&\�\��gM��@���غ:Ud65�j3!*��WG�r�c�K�J���m�czׂ��M���E��᩽{M��k[��޿��	~õ\gW�H�?s�;ƀv�Eo��I�A��BbgY8)�?'*�%���>d��.F=���J�9#�,:����E5N���ܖe}��5�OhۻĨ%�fC�f�LC5��^<idr�R��0���EF����a�X���6���.YO��!d��{�40�=,]$$��C�G�}e���V,����@Y|�+���f�뜛g`� c���i$D��`��:	�C>v�'|�T�+ W����+�p��D?��;�V��C�!/@8'l�&�JQ�We����YwU.�R����;;Y��W�����R��'�ջ1�2_JF/�����c#6F�I�a�X1�]/�>���&��V<tn�����DĲ8c N�gM�R���V�U� ���4�=�;�]�M�$��A8��
����@�/�jfS�.���Mi�9��		�*Z�pkI�>�N7���y��Q:KZ��Db�s��[؛�0O�b�&�����Q� 7T�`h�ca݋/5$�P��캀�q����[�;@F��\I�Sz(���Vr�����R��$��:uS�T�;�%��*EN|��N�$��r�����M��ôG�!k��~x8���-X���<�a�|ps����4�w������׌��	i�����dRuOX�Z�s�1��aX��A��X�Z4��~�V�vQ�.'Y���H��y��8/O#x��Tw�|^@ѭQ�SlS/9�\�Ob)�%;��wQ=��}��?�C�[%X��`nZM��]\vՑ\knQ� �ٙ�'�JUgSC��ڥ��P���{�$J�bi�Oj�����}] �`�����z6Rj�'z��y���c��N�&�-QW�Z�y1jمk*J��*Q�_��� ����'j�R��%9����5Q=�ʘPV�+�vm�P���q��	��;������V�( ��Sc��H1�����^-֌螁}l��ͭ��5.�>&��NlȮ�EqL��fo�=j���]1����ۘ�q{�oV�um4��t��$uf�jD����D��.f��U/n��3_�1��$}�#��F�&�����tU��Y��أaA���ou>jo ��'ᳰ�f�vǮU��*L��"⒍�'Ȏ_�	�4��i޹�2iCh�X�Y�[.>��Z`�O��?1�����_I��T'<�(/�z����s��e�K�Ga&���<����k5�v� oS;�'�����D�OT���$U-nU{MC.�X#)N��������Y�C�ɯ)8v����S;���� �+/Q���ι�z�����Cy�̱w�2�������Z��iT9���z١fAL4o�G8@�g�t9v�;�/p�Z@$:�h�y]��Y���N3�bKO��S(����0'�庄�5�K�x#̆�xmP�dAcxW,�̲�z��U��ÿ��"��Ϟ�k��UC��V.u�\^����� ����Y�?�R��Y��x�[Wo�vG�����}���}�s(�7��!u޻����&F��Y�^�K�ԨˤS���oƥh=�{�)��>G���Ֆ�<�ب���ٻ��'	����*,���f:��8�a&L��gd��]���Mn����u5:mJ]F�fg(�|�>�O+��1r�$�Ec308�J������/|t�n�`аxj��Zy�d���Ȱ$ n������[R��c�ՁI��ȑ��!7�6_��4�/���`f@!�Y�	1��Tz��胩 �W�"�2�E�}2�h:��<���&}$A��7P�;����4>p������߷��_���"mc�h"d��Jv�X����	H�� NNA�O�ˠ��1��ù+G��+Pt�rl+��S�3�I�6���K&iRݦ�ݕ�Y�s�y�.���}�]�	���zK�>=��C�i��gj�3X\`�Kh�	0�M#}�����2+����u�"͔�����-9@|��K�-P9��|̺���ʀb��$E��e�@� �A��'l�LҪZ���aƧhU� o��'�fM\����6�'��ܟ�g��ͅ(�6)ڵ�y�p�!�y��B�×q����R6G�!D����;�~ɖ���]���@����2��h!����B�&C�L+n�D�`#�(�#�.�� O >�Z�x���adJ8c�F&����!�M��_��"d��Ԣu�$_�9��|��h�bY�o����-"���H��7u�>f�'pct{���"�J������]��6���x� uc�X<��~��yj�@�.Km_ )��a1�s����J�Ql'#��s�qݽ<Dz�x�{`�
�n�5J鼯���=�	*�p����m�Kݪ᙭}$���Q�hq����7��q�*3+=��G�X�ᣭF- �!e���-�w&j1炧r_�U��t�Fύ�����'�NE~IL7zp@EC�3R�gxhu$��X�v�$K\:��A��K��{*�c_��EȖ���2Q��~���[������0�yz#�G1�5kQ�����Y�e��rU��:g�pO?ɐ�T��l�r�N%���e��	x��6Ξ���g��jL����[ɴ�ܒ;�|��C<�ZI��&���f����^&<�i�\�J84�إ�?�S�����U0����þK��|���CM!������=���2��=�b�@�ӯ�i\~w��D����R�ޫ�d���4��T%�i��`�Da$5���*�0���|�i�]d���ऩ���Hh��s���u��AP�<��$$߇�M8�6?�~<-��Z͎�޺���g��1�+��;�]:+�s|���s��� J*��K
h�c�A��3H��qi��'�������Ͽ����u~�t���V/�_b�*D=�|�6��߳3^!���2Ə6��xΗ}q���\��چ�	�%�ҙ:��htQ�0Nw���|,����D��J������JP��' Ӟ1�Y	Kv}��e+���_0�<Pj�5�鏵Y2�
����͔0��=�F���)���:�[&͟Z�d5���_�S��fE�o])'��J�����k�/k��=Ǧ��ݝK5ɻ��m��N�C4^ڜ��x}r{����M&R�|���+�!	��(�(n�!�S�d��b���5��
J�}��LY�^��@�g1��ϗėyU�;�T�d��#|�� *�"�ϝ��QV�A�W<�?�b��U�� +y�JRdZ*�)8����_��ː��b�҉���SG�G��8u" &�^Ť����}ҵD�w�=>�璹�`c�|T������ |���ݛcn�#U���2�q��m��P"9���z��߻!���&ʫ[P�����!��E�s˪{-�⃍#�$b��shC��pk�I�>���� Sp����1��0�;�1|2�2��@���!�x�ۜBO!�@eH�x[
x����z���q����+����f���C���t6Y�?<��G^��^���q�J��72"�73�@뵉�55��o�5�L�ϡ��"u�z���!#�e})<��vN���m<�mG�ߏ'y2���=*J"�Tf+ҫ�N�j�j�,�w�Ih*:�(�Uh,{���;d	�.����[�`a�k�qL���(��?(����f�%U���(�ƻ2�lcزG�n��Q�7�L��ZrS�k1%��;�zRr׷���o��w�P7L���U��(���n;*��&L	"r��b�$��N��2�[�ycQ%�����6�28�~��R;��5\+�Yf}�TU�JY�3�wY	(ܛN������W�(Fr���L)��S(�GZ�w�AP�Ac�"9[q_�⹃&a���K]C���J=��vIY����-��xG2&�TT <·���/D��u�+��৑����r�f�2�'�⯜r6|%��9�p`�Ï����O/kn�D���_�ZSXߎ]�tL7�p��l\(9�t��'�TVȥu���I+����V0���0��1�������j	|HaB"
$��0l9�	e�Q(N&O@S!
�F���S�ɛ���Zv2=���voo�r*�B����d}8����D^:�U�^�2Vj�ly���q�%K��ݲ�.d�i�à+�C0����B��[��<�W�ߨ��{ʟ(^'���tM�:������0�v���S�Z�i�6F�񤯖&�J�e���U.*��5��S9b2��=���ն��~X���4������;��'��c`�`H�R4@!6"��)�Z����
`� �>C�~���K�_����G����Y\��Cs��٫�̑��`��\@_�kwC���!�[����Ulc'.Qp�9��\:s�;]��~��Y{YMs#A6�nQTS9�zu��NZuTOBJN>���l�ڠ!Du0'��4(YQ�6���e���fM�W>��!��� ~9T7�P&=�t�܊��<�����i��^���&���B�5���	�U�&^��3���!ڬ�B7���\͓�,:(瘹OV�^��{>:E���G���:�"g!2u��7���J������M@���ǧ���ԗU�v<WyCNy�? ��>�\.v*�R'�\�[+;��%`PXH��bNNv@��P��-:^�*'�f�v�m/�ݳ�)��XS��Ni~f��1��(�O���1��q�y����?����^q�N���5����\v(�#*�SIj�ؗbԴ�KHR,D'i1���ow�D�)q2�wH'���ѝ��5����r�/L09�CSc5���x����I�Bpq�@D�*����pvW �5
q�q ��G�%�'���)��c��]������l*�=�q�Qг�q�����E��
�W9��k���
��[[��<��|��'�n�]�)3y��_�iʴvj�$�ycrE5�>(ihv��FQm"!�����.L���ڤO�� ���`pH��P�(����{U@f�'�0UU�sx�ڷ���S�
�T���?�_�w%K�Y{��1h�EBFl���=ܗo��ݪ�\�a��KumPi���3����>Q�ϑjX����ap�/"B����7&��ʆ��l�1`P^�,���� s�.fB5%�ۜ�`)Am3��*��*0�����HIXMvL�� �x8J��=�:I��Մ�X�y��`� ��q��c��fpC(!Mwx��Hv��>��A�ki���^�H�O+����:(��;�����:�;ȑś�M1�F�[��!t{�m6��ק�}y�*�,08��	0ˆ�y���
�3�tyPߓ��2%I��G��\�2���	\��'�&Ve|I��Ea��ZB��_nŧ1#�Шs�I�`"��oo�fWZ�k�vG&��dLl�'��ObtC��q2��ú�}���g�h̭�lTAf�'�Ud>d���"������
H䂬1�YuCV<���dQ2Ҫb�9-��:�q�w-E�X�Ws��Qg�N��i�vv*�e��ڱ��H9�t�70;���Tv���q��ɻ�!���X�G�'n����.Cq0����.3	���S*%2��d*�'��f	��@8/ZgL?X�g�gz ���T���y�ع�VCw6����'���,�D�+PU�o�˖��A�{RnM"���(˙	�r!у?Y��FR㛝3(w_1zi=!���Yv��:&aM@���bøe��1�*�?l?^��ؾ��:��Ӓf���f@��=� P*�L����|Q���9lu|��f7t.	fGK�L8�᎚a����8�&��;�6�6��K�]$�Gb��j���` ۧ�d��ȏ��$�
�:���ƹ���a=��*��C_� zV����e����<�4������8_!�����ھ��x�[!�˽�������d^w����k�U׾��hR���7�� xx3�9#`��7�a�ڹ�i�gK�'�7�S4����Lnt��o��?'�?�l�oc��4�e7(Q�|��&X�Nz�$ti�1��ǋW��<�Tpv����CO���I��*x��*{LvM��Q��\Ts�İ���=��Om-�������=������9�K���.ԙ���%�%�`&	��8��ٰ�
]8$�4f=��A��y�O���G7���0���@Lk��B���0��P�)Lҷ�ы�3pd�/m��z&��gf���\�D�Ѓ<������#},�Z��y`����,��/��J��#;V����kA���@�E_���M�VF(�������~\�&^0���Hh4b�"�s���T�"��83˃ǎ/E����ˈ)A���~f쎇�K霡Z�e~Y_f耗�諯u�KV�Ȗ�[ͫ���*�1W�XW����u1�]���$K\������c��iD��t�|��D<Z�4�x|����@�!5k��n� "0}p4�лhU�[N=j�p�[��gCH�t���r�x�K�0Bl��h�VeP�ҟDiz�ah��>��i�����z<p�E�}JN�:y�i��D�iԆrM��-���)�����sI�����~��Q��8��Fچ�ι�q��y�����^Q���	p	�'w�!����=��^:��/X�gKS�ea�"�3w����&Bf9�hE�j���k�d8��r#(%����QY�,�]� �.\��f�g���m��
���3��́�%��>���z��f9���F�K	�"��15��#��l��r6�}&����� 