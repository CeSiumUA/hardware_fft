��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�	?G�I ���&r���r�,	7=���b�ĝ�#�*�aØ��ο�H�x/�-�R�o5���u�6%�~����kq��yW�9i�ф���rH� �����|"�9	U#�'�iͿ`,�,]7���0��pd�n�@x@GtQ�����a��o{���'��Z�3��m��i��G�f{n�Rڍ0��3@Թ{���tt�<V��|C��!�'�/"��ؾ�j�X*�#�;���A}_��1�2OjV�:��kH�E�W� 3f�;5��	pR���
&�:�Li��<�v��{�A���!��;��B��M"66FuN�|{b�D�I��t+�!	'E5��mL�*���< ɉ�����`7^
%�
���X�(���tՆܠ+��01l�[Ulr
���S�S���P�65 � �B���������9���<^T��#d��(39������/R��n��
��_}��V��(�.�^�&���ѓA%'R	�~�a2����������7k��t��-���ea�\Xw�	=��΃��X�u��@]q����B�����\���v��s��k�
��ůQ§��"lz���Y>P�Y�򯩘�u���IzT���Ž{�{��h3�GpoTZ7��\���0�ƣN�u�>,I���������0Eht��}f����?�T���b����=�#C88�)\`Bu�%%�o&(:���,g��[�I��>���QU��z�g��X��Gw�}f�r�-�^��=Qܮ�X��4m�_���U^���=�(����W�=�=��L��<�M7'�tL�|ſ��ʹ�߬e�5���Ĳ�����7>�Py2��˄4��3td���.�Jh��),\*���"�k�S��﨧��X���坴��({+�S�\�y��[l�44��N�q�Oę	q;�$I5�TL(�&��f�ħ�f~�����Wf� ��?��L�$Օp��䂠�`H��c����3��e�L
F�N���r��%��Ϫo����|n�yQCe��!�Ġ�)������̸{W��ϭ�g������Rf�[@/b"[���`C.@ڜע5�-�@�	uB}�`�~���>�<��&W�oӚ���N����j��]���58��h&ۜ,�L��q�/�h�{����Xz�6e��B0<���	��>�Z�o� b�eω�H�?��~�T���f����>rm"1V���lE7�{1䖉^{1m����6����3�����D��A
Ĩ���c���?��Ԁ��J�����6-v�͊�/��3x��7��6v�r��D'O�EKW,σ��/���	e�)���\7�=\�}�;D�<��鄐Y���de��3%H�ϣ}%R�BAW;�4?Nw�w�V�83{p�_ VH�F�U� y�;�����_uŧ*�Ft���%}r�5��J�i1YޢN�F.	��8P���?dTK�;]�x��(؜A�;�N���&N���]�.�x�{U�\"֒>@�KX��ޱ]%y��@��*�z��&I H���uY'�Ԋk�lb���a���Ry$q%ppЙ��Bbd��D;n-��=��	mbmP��O:QN�����H�O�*�F�[�u1	z4�9�<8��+���q/c~�Ԍί<DqC��E�B��)J���kf�<���/�]����v�AR�� a�,�j��\,�y�T�OWNdG�A�v_�5�LB_�Ǚ��T`���*�Gv����n�%��G�'��QV	�-��~6��E�0�Q��G)+r�S�V���\�5W�\���,�E�B� �#��5 �5�3NY�G~|���Gn2-tVzk�T��(Ȝ��=���1J2Y<�z�#,��㵍�қf3�ݽ%ּ3 �aW�ّ�N������{�?i5C��;�3�05��\z=�.Wo��� �(�sD��ݤ�f���'#}�*���wq���IV�Պ��[��s�O���5����Yp�1F�{��3g	�"P�\�ԛ��[�h���*����εiU��XH<�1!��`��q߀S;uD���k���ڰ���������(�d�����n!�j�:f�yN�ձ��5�W�G�Q̕T>H���b�p��rc���(A@��9x���L	���]ٜ���اd[d�|����dK?�[WaJ�	*ݦ����G*o�Mwn_V�����$�i�T�5O��g�S�\g:��#���| .�݃��
N���eQ�,��R��Τ(;/��7iU�i�X9�K��C��:� ���a�|>�j�$����*�V<<�jd�� �������S��i�ʰb�;�Tk꩘�S��}x<�s�����d ���0��^�tk�k[����R�06����Ώ 櫅=�ѽܻ)nyB�f2�`߬��E��l�6aupQAN� �-(�RN2,���+Ʃ�3#0&�v����i&9�vҞ["=i�;@�UO��ڨ�1����Z|7��d٤�U[\�IМCoބ��B`�i'�l���]�:v; M�����L�$�Ju�$*�����J���:�����r���<D�_����]0o#�B�+����&:8EJw�)��~�.]'�Ww��ܳ�b��IO0d��^�g�.d͆��h���w�/��謪Js����,	K�$_o�;��ք���:�ײz�E'Z��`-��ſ!|4����z%��5b�9��+���DSr S[��R"�HXn(��6(�Wc�HL�� �� ڂ��]���o���pJ}�`�=���Z��Ղӗ����1Q!W#?��<o
���	tgF��6����ƚ{��d^���@�
����S%���D0�x7��ܕ��j.��]N@�6��# ��U��'�qĐ�Mog��.��t�:�
᤹���,����	�K�h�Q��,�!}���Eņ��}��/�2��-��ȱ%E��]�|�������T������T9[���o0!���}M�~Sr�2�^e����[ƀ�"�6�CK��p�<��nBJϙ`�d�,ԭ�,��̈́q�t�$G�����,z$Iq��MMm�Op����b3 �{\�v��/��#�$�v
�k&$u��o��Zb,�cM���+w��uK�S�F>|�C����B�����S� pe�7W���,��Pnti��aXO���X��,�XA񜟮"M�)BB��A��e�%�������eHċ�Ny�i3��6r���4Hzk�� 7vZ���jJ�S�(0Ĵ"�l iqZ+�.�i��@;�X,~�-�Aч��.8���GZ�'ŵ9��!W�s񚼞!-
D���3;� D�aX�����)�u��n��յ=f��������9����<k��W�̥ɯ�O�[h�r%cS���K���-dEB�Y��S��ݼԯ7j�������.���ހM��LM��BW������mW������4��$�RN��'�dTy|!�r�ZA���?�( QXpN&����Ey���J�s=Eۿ
|K-ʯρ]��n��x�\����
����k��}3�$&�#�b�c.W� 2jݣ�<�Y�͸���a�{
��.p�)=�p��F��$n���N9���� ,�i9�ۻ��d�c�7�]Ò/�:�Z>�G߼_n����JsV��R��nq`�LI�i��L*a#���^<�l L�
Ea�pͳ�zJ6��_u���x�~�o�H�p��߫�����`DB�W�]���]1�5ZICQ�x���j$���"&�C���9�V�N�ZS-�p#I ��RJxe���#V{�[s�TA3�����e��a�o���Ǌ>"1�� �7?��بw���9,1-'��)@���k�_��4�F.�#�u0�\!��o(��G�cJ���&��)�G�MLb��S&d��o��5��f�,�w����F_t}�V܉u0��Bbp�M/��я	<;�r-jeZ����5K��ꥦ3��G``����
�ޠD6l�`3ɪ5�l���u%W�bH�.���Q�?O̙7�l۪�\���D$�x.���xN�p�!Ռ4`JG܏��������a���}�K������uR7�Kqv�JP��A>o��/��z�W)���������#���?5;��XLﰩ��Y0�;�hO�4i`Ix:�o�]/���g�I�B�Z��?J���ˈr�PRS�,���)�sh���xz^��[m^�w���%7���p�;6���$vs��2�耕p@Ȏ]��YC=Y����Q-:�vg�Id*s��ߛ}��ڜ@�<����
�A�d��W8S �A+x�
�Y�,�r<�Q�F�(Ix�ny#w�4(���bt����5wI��"VZV��kԛ$�UM�fR��:�v�^�ۡ�R�CX�4�s�n�Y�2���iaB�n����Oh'���[F`�x���P��f=ip �U�㶿1���T��)�XR:�>�y��yLXv���������%���\F��&�6����TiL��R�EM�}��1ΰ��z�˓\3o����q˚w�g���q�:&k㌲?{i��=B��R3��(�a/���?:U��*g��[���P�e��M�:����d㶐���m����J��{u��P�Q��
�W60�Fp�ܲ����ĭD�`��*tt�<�#����ed*�G�e����+(T����r̕/��xi?����r�(�x��X���~�H2�Ig��qn��Bͼ��������j>���"5 e�`o%�p^m�%������̵A\����h��}�5��i(���g"�DL輥۔h�¨O��(�Rf\t�[����4p� ,��8y�� 0�IB �4���̾�wB.��_1<��!jS�ֆr^L�5�˭=��b1vܕ�U��:Y��.���S�#��9箮u��Pc��	͍�{�0�*��i�Z��U<=MsDl��'Y�:4)�������l���+/�X��ξ��H���RDG�2��Jq�E%R�1듺KXm�_�,Q�H����ker�m� ��_ɫL!��$�m*��R�H� mi9$����w7�E�6��� %#�������o�t�ܙ�����\S�
E"/�!��E�dr��p[�[ŷ�|��6�p����fWk��=
y� �g*j�e���*��2����l�4�63x
�OȾ�t7x�A�������`M����AP0b�e*͓\M�����4$��3�v�%0(ʲ��{ O�{���?�lJv� ]� �FrB�t[h�L�@��!.��9�3�"-�Q;��6�P����r�ϩ�˳�$�a���К΁G2I;�o	�t��\؟��`B� .;�����(n��%��xCn���M݇�ᅻ���5��,l���XipGK�Q�EC���D@�ɚI�{�$�c��%�e<���ޮǪ!���qꝯ~D+@ST&���?� o��,L��..�d�/Q�2��"���[@u�I
����:K�[&� �j�nqx��3|�&X��mI��ҪB��N�9b7�M����Kn���b�zNM����{^^���#yb��b0Ot�#��a��u�gR�ل	�]A�I7-"�`�|^/d��S~�Q��\G�>��Ӿ��"w�<P��Q�������C[��;�.�Q;*�.�b�W&�gPf��7�]E��P*�XGu�oQ�{up)-@��7v5C#H�v��Y�R�Y���)��.P)�o`���ٝ�(����AP�ݳv9��ğ���-�Y{��[S�34PgĜ�:\��|sd�?Q	���,���{�D%VB:�oZ�>Sa�5�g�dC	�ܨ3^F:���٦�ӉDoE��^���˼�͐���)��1��V�+-��0a�f9�ED�j;{aף�A/�pi��_@,S ��=��O4�������47Д��^#ܴ!�Ӽ�\`{�r;WwAW�ژ[�Ώ�3��wƘ<�W�����a��oum����#ﴅ�L��̫�<���{�m��~n�����e��(� �g�l�ѷU	�ݗ�h��Q0z@L$�T��bK��:f������;�y.��B(�4�g��{3qS[�:����\&޳���'��-0(L� +���õ�+�|gL�O����߂�������5�}Ʒ@��Pl�����X�̿ʙ%0�{s�=�8Z�c�:��ۍ�(p[z�ѓ9�Ei��K	��Z�༃���a��Z~)k�N���-*�lϭtzmM�Q��D����b��V']\Z̷Ҥ��oj��+��<j�S�{=�~�?���kV����L�e���j?���Ͱ�@�w%���_��5�a�IL������X|C=��|����4�<�ŵ����N
C��i<�b������n4ϫ�|h�SX�q��˩A.<�g��ؾn�V�0d��)yt�S�>U��*���ٸhxc�T��1�NO.C��%j�����=Tj���9�񳡴4�DbM�)���r(H	6{��R��c����"��/k��_��W���:=��uR�9)�Y��Qɤ��XT�M�1=��%!-��`�(��s��ic�ü��͡��-xC�w�>���S,��������F��{
m�ݙ:���� ��)TэDf�\:�W�pk�],��5�r��������z�	�.�V%踥�| ��n�j�n4қ�O����v�=b�(�^K^��t���Ɔ��󀖔��6�����I�������~Ǻ3v���52�,e���� 1ÖCu*@����E%!q�x��b�����H���7�Gm�|)t��7_	�ݛ�Vce̫>��z�y�W2���#%���WݮfE���l�m�1.+��2��'ZS�����CZO�GơMU�(t���Ȣq3�8�K�m�y	FY�+����97�fD��3��u�߻_^�ě2�Cg������ֽ�ؐ�w��}m��d��;����w)�v9����9��Up��+�|�떬/	P4{!���-���֒3���u�R��Ӱp�k�l�^+����@�$�/�b�z�ju��5o�yIbFC��ic����z�RQZ��)��"��f�ŝ~���$��=O ��q��j\���PRj��VTC��G��̌+¦:U�>�˶'����� ����w���2|�Ņ�^Kd�o����v*vHΙ�7��)������y��y�R����Z}��Ƚ��]�5b�($(��� ���q- ?t�^�ȗ@C
%� �X=�����bSH��K�L"&f��=��E�f\��,�,u����lXYc��a���^yA6�t���Rٹ�~K�	|�1���z�3�ܷ4#�Ur<�ӟ"�d(j�"�Px���mq�w���IcA"�kSp(�� "�m�jS��?�a�/�[2֌�+k�0R$�׋œ���W &1[ft�w��9j�aL]�%��4���F�4����\�`�E��4ubr�ϐba2z~U ��P�3�:�e)C
 N��{�o �|q||E	����r��C�2��i7[^���R�9S��p�m)�3��B�?��kƌi��S�Os�t�_ט�9L+O���v���[cGw�g��3��TS.e�r�7�r�/y&6�5�ӥ�!�j-��Q:��l�����XA��`7L�i�"vۀv�v��H1b��0�vސz^F���&���%�  �U�hVN�F���]NT�E����e\+�y|�z`��H�U�����R�	À�����=C`/�1m�p���F4S�L=�?Ӡ���ol��wv����|?��2~�ۛ�IU���0,�Y� 垻��1�5M��ʒ�}'�E\���DR��K�`���_���L���!R��l����uW��ZZ�I)c!�چ|Kgc�k��7rH �eq.�3���릪F8_GŊ!:�K9Vf=X�0귡5��n��[�{����{I�PB{�HAU� |�/�O�Ȋ�Q�G�̉��^��ՇM �A�'H�J�U{]�%+~iM�����K�Gm	��[blt{��no���/�ݎȖ�j�kS��	%勜ҥ��ԅ�Y����>&5�&��Ov���Ni�7HH)&*m��^^���[�\�x����-��&��75@�\g��b���ND��l(�W�/$V��i9c7�Y���.��A߈�9�j��$(�'��R%�*X�"�=è��" Ӱ�}Z�?�k�볧��i��px)@�A-@,\~cC.������*dE�ٰ�����4e/�抓bD黿������+�P/���#��gU7�8�Ź����t(����BF�8���D+xw�ٌy��%�O�+��	4p$�}�ʇ�l0w��Pқ�-}a)�%�uZy�_c���==�\	�X��Aҹ l`�nɀz3xϣ���@nE>���G)�B��i���Ux�8�c�=qQ�i�� ���Lw��ߏ�މ�w��^{i�T�m�%����/m�������疕*�ڒe�NS,j�$~�\��T`�����;w�,T��1v@�v���h���g��H-�&Z��lz�^W\�T��s|ɸ��e�����ԝX�W�vHK�~,�1�<:S�򮁓�P�o.jiF���Af��	�)���,�s����J�ai�s��ǒ�T��!�*��	B�2��$���jJ�p��R�nM�ܓ?�r*�
��n���j.)��$Y4�����m�/�a��Up̠�T澾���h��b�r��V��C�8�w���Զ=��	h�h� �	D��Z�W�@��;�/�j��W��-sebc���O׏;V�B�B�ӥsFY�.H:�wѷ�z�q�#ܧ�s��NN6:.ـ��Pe'�2��M�L�7�ݞ�Փ�C�^�)�S�v����y|������d(����߿=#�*}pI!�C&����*
�C6^�[�!tΛ-�#���M����K�h���3lv9�'A�8ز	� ��m� ����{�Z�� ��&!�}T.�О�i�?2j���
d�&XT�z�=����Ҧ�}��0�)s?y?�r�^�P���i�qU�R�F�q�����"1vr7���!l�8毰H�z��J�r�����i�3�C�̆����,n����*��t&F�D\[s�w�k]�Ӧ��5<9J#�|��ji��<��K���Dt9��^�ǿ�(� q��[�0zm
!�HN[u��z�m�QU��#@��q=��B�J�I��3���x�����Ƿo�ļ���!M�8��X��?�Rz�8�x�pe���9��*ff��e�m�L~1�:��,
��0agV�ȧ0�{H�Ǥ=;/k��y�K ���׶Rw�ݦ�bV
ɟ���jl�^&�8����FEˀ���>� ������W���+	�1��E�|� ʠ�3Lw����6����CxT$	���e� �d.�; ���ُ���n����>.!j����B�zL�`�pr���"4V�8=��O�?͒^��cCe�i�S��I1K�]R�{N��7���āPo�Yf$��z�Ѓ�f��ʬ���+�
.�����H �X(�@pqۭ&�p/�f�����X�o�K+�Z�O�P��������O�<wN���B+�9V,�6"U`�In�a��Ć��A��k��~-\�����,*V	&t�%K=g7�xT�$�Þ�i��-ݭ|"�|���pg��O�9��xF�����1g\Rfɮ��6���B	h�
nV� 냝ar����q�/c��Ƀ���i ���f��?R�kk"U_-�CK[ك���x���dj�·q ��O>Uﱁ�B93X���3��'4����ڿK���G��Ԫ��6�9�>V�q�!��	�X�Xzk�iR͹z�܅CA�}��"�j}�*@`�p��B���^e`\��G�����ғ�Q�z`�����[�B{{X2�#F�Q���~E뚃X�!�Xt)i��īM�bV��g�����x�1tYڝ�l������	m��m+�w���"f�\���鍮y�i��ӡ�;���X�6��� 3$����\�$&�o��Y<#���t<��(Ug4��w�� ]�E^�x��h[$�Nїe;�8�U��3:X��ެ�?-��qy�x����I%Uz�$�[zBTq�T1��v�8���2��X���z<f/��;w���{��S1������3+��U�6?��R�V�o}T؃CP���o���h�r�� �mf^ĿA���T��j��q����n/KD�fͫH����i5��ix�����t^�l���4��d7]��%���b<��B��@��jfq��@oi���O����k�G@�L�u����zP3�����(�e�?ǘMtp�ó��<�q��ybUx;>e��xgx�Ziq�bMO�����2�WS�|��Wt��=�7C�fg:�W
>r(p�*t����MW�aA<z���x�Nm:�I3�݇��w�>P��w�U#2S��h����v� ;�gL*�n��]\蟏���K|3��a�Y*�� T-lP�[B�K'�F��q-��7�5�>��R;�YK2��x�Z�:� ���� 6��AKK���-��Q���8��r���9b���?��ȉ�KA;[�+��g!~7c3t�./e����`1~<��k�]�cz!f�Z� �y�L�U��I]h�}ت��GWX(�>��a�#g�gU-4k�X��{]�c4ݔ�6�����ݠ�D�DF͞��/��!*ԍ��ͩ�����MϹ�Ip"�K�Y��,�`b�����Оt���	wN�`2d5��0�M���|�,���k�Q6��<i�0����))�Ͳ�Z?L����.ޕN },p=���۠G��/-Q�߷�/z��$����5�*S�*��u�N(�p,�����Ը��P��!��O�i&A=��S�P��K@��^ndx��d�'M�{�^���͛��\.�L1��T�G9�GM0�"Ds��7x�rݰD�/��;���+7�[f����_D�i.�_���2^aD�����mm���}=�й���Y�3���
�U;V]�+�l��<膝 \�d>\�fٛ��e<jzCݧ6+��KV���-�X�N�Ҙ��4!����?�����<`�8��{��K�֨�Jw-2E��0��+;��A�Pb���Y�EAh9��n`�}��ҥ�خsݝ�?p�=#����7)j� �uEГ���r])�3�q�Do��cK��􅵼�ʾʺ�-g%x=��X�)�D�L�_��`͈���j�r�E,�+��w�J�K�X����O-n���<lL�x/���,Ĭf��EH�H�d�qA�W��{�i���E��㇯ܗHg��Qѓ�8^�B�p��<_ �A�{���g)fεPfa?��7��0y\�y�z#�M��Y�]�3z�3��>p�C��q�R~�f����>b3 fK%�w����T��5��μ��b[X��񁺲W !���̨�E"����";�I��)��(�1ډ&�<��q���u�r�J��q�Yۤ�#4����D@2I�������.��Ylb�^vO�/9>L �Q��$Pf{�e��CwS	����8i4�a�~?�p��gW��ؔ:wSh/<nݷ93�CD������(V$�۪(�ҋ��Y��2g��ѱ;��f���\��A_�GJ~���L3Yj,�,P�E�/�����8]5�F���͒�j�����:�l-f��ɓ�����W���W4� ]��6f�呆�#��:���2m��@(jK���y�oM+v۷���)�Ǵ�lu/Ġ�.4�T���c���&u]�b̯�^*yJ�m��5z�_�l�����p�m��qH�@�7��s�8[�&R7G�ׯȰ4R wRTu�*����1�C�0�BL��ăa5�ao�����Pz��w�mے�jx��������M��q�T��~���b58`z�Ù��%S��5*��B`�#����f�E�J�B�?��!〥�8\MA�|��3{��(>�Ј,U�&�4�=o@yB����A���'������
�+"6�M�hw���Ê9{��TU64�tg�N��U�k�>��'�r��}b�Ħ_��u�%�{GL9$z�y3���
��!��KQL,�jV.֧����2��%�L�s��p+ Ă�	����
{Ƌܛ��K��/Q^��DUЦ}��:4������BI	�l0>�������s�I�l�ܬ+��k'�*{��O\��h	e��w�3�9�w�z�v��"���������+#�������颔\���������K�B"��L ����P����E��� �6(�ZV�!���wB]�[q���Uyf�#{���E"ӁK�8~���eȗ8���.��ۛH�Z��c�}�D�Ǵ�{��s�_Fz�>�8	�zϷ^��b�9�y�]�:#k�D;�委h�@���0M�a6S��ޘ�� Y5cȚ59�'gMS����P6R>�w՝���	�{6�c�uO!V��G�l�Sx�A���������D����`�B�9,�r��pr��0~*%�������R�c��[^��/�Y!����֓^W����:��(�j��}h��^�i�ex@l�~�L)�9���&�|!��JB]��:}e^�T�B1�(>q��<�}��d�-��_D~�
���b��$	�|���1ű7֢?/h@)����`#���/��1��-��X-�.��P�d�n)=_�T	���.Z{����_Y��kb���>�d@�4��7vV6����
��	9�c�[�v�<��]�u`-Yv���� ��v0M��z�� ���81$ʤ˩<�����6Ih2�r���3-�^��laJ$i�SI,#�ti�?�\y#J�6��iwm�X�K<b�ebަ�w���X�*���jG��eӾ��K'�̿ ����]V�iz �'��A��|XF{�B��R���:U<��3��u��e��oˇ�Z�L�g>�D�ڛ�E���}~j�(m�jY�BZ��Q6��-�e��Q�ܞ��ɮY�tB	e��Lܭy�:ًP�ͷ�]ۥ���Ρ̼�e��u����1=�;�/y�7��t�dOM^ݙh��9W�;2ٶp;ȡڻ�y[l�"��Dds"%Z ۞��Y���C�
_|P�5��Ѡ��� fw���I��9*����3����{X�Wm:}i����(F���p��U�P_�x�h�O��[l?M�G�T���~ݐ�������ɑ��6��,�xm��F�V�6_�i���ۜF��t�+�W�͓O"�\wZ�Ig'A��N�>lq���,!zPL쾙�.���+X~��[�?�n���z��;uO^��w���I������=2��D�#��z�o�>)���U��T�^I��;�bG�$���N ~��m�Z���N�w%��cD��ג�BØ:���#5�&DZ����\�z#��M}B�ɥ�[��Ώ���vs?�v�{>�F�SÝ)�gq�K{���[W�q��E������6�X�W�m�/�@�x8S�����+��	NI4����7��B��W��vӿDZ6��
�j��|�Q��/U,Ǐ��j�n�X�2Oڻ0���LJT�l&��`����h���
H��%�����B�TB�>z��.��=�W����Z�~�d%��)JO����MDʧ��ݞ�y��(��s$0��cM���(n����#�ʐa�~.�o�ٍ�Q�k"�wR��mp�{M�~J��u��3:/
�w�vD�W�7�̨���M?y[aXtc�~�N��n����(�B����9sj)!o�&u��%�6&���Ö��,���zp�k����Մ������f�Juo�2�n�w�R�(�s�� ��E-ᘾ]gkWP�w���j~�#(!�vr�����PC� Y�p�D��L�-�ټj 0m�"�jd��ݍE``�5�S�`�x_d[F��ٿ�-rW.�%�_�D������\|[=33,�bz��c��N���,���얌"˟�dM��h��o�q H�^�j�*d�0�cc���,����/�w"�ߔ&��9�Ü<�ӔǱ�������#U�&!�ER��z�H>�>��b�k/��f��B����L{r$����l���рM����}M!��%��AӐUv���3iǌ-qrwᜪc�S.�V�>�{�����ձ+�lr�y��������(�����C��	R����7���]���M# ��iɀ��՞���@�{���U2�9�6����Q�tr�D�C���[��m=� G�g���Lc��v{r��o�B��g&8H��W	(�x���'�é	�i9�G�I;�=��)�)W���ʬ]̋�yy7�~�z{�Y��(��#"����ٞpS�-�Rq�ҝ!��Dx�4���l*��+��T�9�s)�zu�T ���BSҾ�"+x=`��y��7TF�a^�|5>W51�{�����迸!��a�q��`�UyP�)hx�����H:�ʆ����k{�&�����ڪ���D��t�&#�3`��l���×�rj���(:u��8�y�\NZ	ސ _��i����$]�m4�@mI��R��@2B__*�2�L=ˋ�7�����F��ћ��J�Lލ�D�M����SiDL��l���"���luf���wg>Ϡ���bnUad��4l���Тi)�)D�w�����x�a�`&5)����OĢ<#)=�%���:��0Е́����&���Ce�Pn2��-X�!TE=���v�_�<Kw�"��;	ˈ�E���i�I6|X�᥇�fw�v��u���2������ S�!J4��$D�+�N,
�^9Q�k媤]��`=dh=��v\�]�:�6��Z�/I�5�*��"�B|~<���}y)Qۮ�NE��{ȅ��~˙���J ���gd�i?���V����zش0���T�>��t��E�����&N
�A�>�Ez�Y*�C�W�l�q�h�a)h�;�܋h�@Y�DA��#�3䜡g�.��}�Lo+!�<1�|��0E��F�J��`(U�>�{콡0�F<73��.��j,���po�sbq���|Îq�Á���O/�{uxW0��-���_�b�;=�e����VΚ�,�6�\۬x0�
���_"V��F�n�Ұ
�%���!#�BCw���ppE�(lƞ�p�[O�c&L�­��RT+v{HG��ޱ� !]j%�H��>�f��<y�:�'�6|��tm�0�B�r�?��9fX�v�M�(IP%���W[1��j�
�,̺��u�f������IҮ�	>6�y�i�m�9�̝צ��cd�G'C�A�ɻ���ks���B	!x����mH��z���
6Vnr->��i,��<K^)�x��Ho���E'����(�0o�Q��n��0e���%�?��U�]�HF�n4�x�3�Z2�qxUj�����b>���^��r����[#?�P�r��4"�.�Ǩ<$rBR���[c���:D��m�'��]�'j' R�_ק�υ��LF�`]�{�M�mLEx�PXoVtZ|��'֤���j(�eh�7 f!��� L֓.V��Q�#�*�9�ާ�#����Ҭ���Wb�)���b�f��c{P_tv�)��Җ�!�#��G�����Ҵ�����Ȉ�>A4�x�!�,��2�B�M��GF�2��is������K�G|�΃�_�	B,Q�^��6^��No/(J��5�U�����1'�j=����\��� d�4��f>H���-�yV'H���R,(p�A�-6�W��Y��c��� 2�7���)H�ŁeU���B��'�A>��, )�ά����q�w��3j����\i|%K�m�ܫW7�'�>�b. A���Qf��O}�3L3X3"	��?�	��R��d���N|c_�=��]����}�&,���8�H�E=ق�WDc'uW��:�Ŵ@��.��t��P��ԩ��>ڼɖ+��賊�F1�Z�X|���^���TZ�(@��;�m�a!�1��Gj�佑�u�RM��8���}�U$A|��{Z��3Z5��Dz�C�Q�^���5�Kx���n�BzU�?���`�h	�K��"�kB{�%���:����{6��SEn������wEtON��^�ǩtm��Ze��]�#�z��(
�$}���D4���o�gc`a�e�L���d'�)I�;�m��}U;�:�E+�rr�I�$w�&�?��A(�Ɠ6:��OSsH-�$����|~�M�0�����a���p��G��S�����ߚ�'J�.a+N���D�Ʋש��H�����"���~0?��;d��5��c�c\[s�Z\�>ì���U�2��j����~E�\+��0�p��ί�\e�z|[}��"xX���C=�xp`9�����RW�X�����+����yB(�d|_�ߺ�[��%KvݘT��� qy%H�7���(���3y�z�Sx����壡�X��;�ۥĝ�ùM�f�'!����z���v��������_�iK �/*���J�Y��49B2��s\�kaw�_5��,�����FD���7�G/��#��2�"(9��g�@H��ki�ֲ{�ߴ�@�|o�΢ Xb?���.Ȍ�Y����F�e؏i�p���1���J�^]d��;"�-�6Re�bJ�n��Ɂv	jJ�xl;����
�WSC��k��4t����a$�~;�槦GvB3k��.r�'|Sc� N�=/��J����r�?-� ��I��PnI��+&%#1�F2���a�������O�jUQU��C���%㎯��4�t��f$`s<���L2�G/�f�37��/�D�g��7�R�����JnW�p�<���6YĜ,�`�>Ñ�0^�8�B�>.T�H�Cm<	��P���Em"�0\�x�;e	?~0v�f?�$�SX9��������(Q���Dਜ਼���h�D�lY���yO��y.�U�>��Ħ�!솧��%(�ӟ,ˠ���MwѱY�y��u9.��w�.M/��x����\��J���׌�U���5CC{Ջ�NFJX�[oK���l�8��,M�̕;pj�����-m���-3&Py�97r�_�L&����G᮹
g0\��M�tZL�%V���\�v�'VO*���ĂG����n݇�}�����S� Qϩ���S޵tT�\�}&Vd�
`}v��Er��-�����N~]PG� 7
������KF�j�����>�1	'Gч�'�"�s�#š��Eswr��1��vv��A�c�g��tq��2z��ʋb�O��W�!�S&�� 
Fh��!��!���g��h5�R�h˝� �r�O�T�3����k��4�[G��0h��S1�Di�Zsl����L��#:�,�ڃS�?�����8Q�@D`ѧO�����U5m��0�BC�a��?�*B.��R]���VH��ա�Z*�
M�h�Q�y��X��J�o�}��0!�۟�$�<�8'G�삤�����;+M��Y1!B�9E"�C���{�w8�Dn��&�w�8����c6�'����^c��1���!��)
?½_��B%��\i�a���>��ᚴ�7��\�oO첀��:�$<�󺼷8N(k��/�==.�R��� ~�?+��Ys�n�׸P�w0��S�κx�r�[=�uE��?GW���&5`R�60����-������	m�x��� �&ӑKn���)��8��Da�D����i}�^����#�	
kB�����͚	�]��*����S���B�ׁiܘ��nىݑb�ό=i���T��������*8�0���Zm�sC��ݓz,�":��E�*�q�N�:��a�`x{�#�{&���{^�:�q	�P�q}�����Ŷ�X�Sx�	�hıܭ�P'_乄���C���6��7���N��q�=�k�b��a��*8�:?��[�YS����x�����ʫ���q#DpZn�<ʐ��H���H_�?�麷n��\�}A��^�
&\玤;����<e#�>	 iX{J��U�t�4z'//�TMڛע�$,
�ի��q���4��[��q���@�;9�U�s�r%y?�/��vjCR�:;��Ap���tb0FbØ��}�
�-m$O�r����1�0;�/k��I�.�����HH����s*�o����^�s��{�u<�'H`]�L����1-�� ��	Q�?�)�F��]VqL�d���ww�A�?X	���h�ɏ�X�w������-��l������P�L��L��9�cᣬ�(�,�D�o�s벿��$�~y���`("z^�����e�Ǩ*�1��R�^�L\l!��W 8�ooM����T���N{��ZR\��p�z�QӉ�����VL����h���a���&�'Z#�%����Ȳ�o��ݓx��E�P��R�x����������Us�?s/����U3����Jr��C���@<���' �'z�Y����ОJ9{�4ǹ���3� ����
��<ƺ�'J=����ԾK�a{Ô�^z)O�����2���G�-��h���hc��"SYYѣaf����Z�e�O��wAo�?Xb��]1Ư�tw$�_h ���c=�����*����j-�uR������j�Ed�/���V�ϧSc0[��{�6aZI�(9i���*��y-��=�f,�O��邽[@e��>���_���Upe�Fc*$�X.�o5&�=<�_?[��,��%�|@�^�P�`-G�-���Q^���DPZ�a���Y���@��^��L��6�1���������n{��h`��5�����������w�t��Oܭ��@��{?>�{}��C�IΒ�	��uv�<#���b�8�S�e�( N��J�~+k�!
�g��a��o��0��\��t�q��U�S���M���DC�T��o���nq��h�M�)%{�I�Oj@o��W-��ii�E���M��Uo����<Aŏ�:D���D��l&"����;M�AͮBA�5*Ig!
�#�3-5��X�^���R��8�ŒF�a[�y+D�X�����]���q]������C-$%[��Ee��,�;�����=���aƔ�w)r��J^����t��9���P�{4��AT)��O��R?�3�H��[>Ci���7����-��A�S��>�*��2c�dx�t��2`���{�xՂ��r�5�z�7�,���,ۏ!�~k��� o|>p���T+)�׈u=���i�Q������x&�?Q��^5/��e��!9�c����9�Oi��{�}o��zfP_sNAMA���
�F���t��	-h�>8�)o�撍(<�EM�jb�<��kᐫ+8��w���8�;?g���p=/�._�{����fd ���2b�:B��'�Q���j���1"��w�Cq��,�@&Ia-P�҆>��>5�!�g�q[~PwE�Q��}�l"@:���L�=��"
 B�3�9Ն�tA�bV�&Z�{�8F*��||@����1���q>Z�A�i=�So���	*���S�όȀ��R� �^]�2��I7Y.K��+�ł�^R ��f5���˾(<loHpn�6��:\���Bo�5��[�px�E��RE�&�1�������
����mnV8D�eIS���j��F6�����&��$�I^�����0�>q���3�6�UJ.ڽYr�L
}<b��^Z���zs;�*_K0L��>f��M�Ǹ�[h�2���/����H����N [�V{�{M��q+zS܇�e�}���9������j���,;x�4��%VT�Զ���uY<Ir{�j�[�=�۾Զ�+�U?l���7���=ΰ���YƱp �I���Q��o�`@�F=e��3#3ମ 4��������q��z�-���-ĝҡ��� ���������C��(�A#�≆Z�ٶzt坪ql*���OJ��9���~�����)�8I�IaK���|�&��I�zb[��]���<-�%׌��E�&��_���kl÷&o��h�矸rWpe���,>�,�l�6���e�,���ci]�f�>��*��������@CK��_�� ��*<�.K�AдI:�"2�P�N���*o�~�r�禚����g�.r��/����@���jმ,��� ��s�Uл��O@^��H<�Z�̞i:=�=,@�i�������_��8�@xJ�x��GP�2 �g�B�R���#�@��`�l�)ak����Ԫ,�o�O;M��gJ�%�Z��\�м"��.� ]%��4/a���;������5�9�*�K��4�#�@<���H܆It���*���u���װ!�H8����+�?�.���D��?�{��N͍E�"� yD�ua)��æ<�j��y�j5�>���.Xg��g�-�1�/9Ĵ��"}s���S1��h}���ַ�	"��B�F�~��Ї1�0ߡ�aR�o'�Ӧ�
P[X����Q�R�j�M�(���C�CKΆ��n�:��rTSҠk����n�3��c������r�����-&Պ2�2�V�b�n`�лe�O���E�*����vK��Y� �e�A0���Т���?J+Z�/f�7t�m����3�{	�7��5�l��?׷y�	*��:����ao��b�U��e���P�I��ޡ�%4��wx�(������o59���º��/P-���~Q����Lw���Z&c'mTճ��e���ZA)+�u^b|��Z��mFk\E����܄c��(�$�M}Emq�$͉}8�'�~�j�1z�
�ϡ�R��P� ���CJ���ɴk��y��ytQ~�7����2�j~6�m"2C�e��<�uh��q/��nS� ��s�69�%� >?�����/I��Dig[D��|�/ئVh�������L��� �!�:��&�{N��L���7��)�a�3��։7��w��4R������T��@�.O���
�|I����_j�3o��\��8��ק^��q1�GNF
Fñ����G~c��uǄ��$>�玘��LJf���^��|*zė�R�-kVAΥ ����+zƻP�R�?+��<�/���*�z�s�ϟ���7��cS&����hܠ(h�Ԯ4w`@V�JK-���X=(K���Vta�*W���sEe<� �[��&�p������3�b���wX�������4n����8b��劢P�0H<k��8O��ݡ-�����Thkb�isf�\RI<�H��U۾�*�צ�B��V�����U>a0�K�9�!ڪ兤��e��S�#���u��@�L����5�}߭������_�<�׭N �H�^����\ƿ�?��.��N����.!/$+�W[ܴ�Ǡ@vY?Z�C�@�A���"qSD��-�q4��MtL�׊���Z�O\�4X%%B�Zto��2o_n��^B*�ҕB�%��1���+��zC�DBY"�:mB.�I�&ѩ�T�5��{ʓ���J�K���@H�S��y#��U�+��`�y7$E.]�Z�@�dc)]��)��b��衿��Ǜ=Q�~�a��:/���շ�"	�ׁYbOe�*��C5WIUF�N��m�;���^{2�e�?i=�L5X�п�����h�"����ڼ��A޸�3����Ip 2>W��3�۸jgJc�$�<Y�ۇ٬˶�Є�0v����Ff`vZ���0�_E��X�	�C=g��h ��v���hl.=Ii��w���c/���:ϑ	��Ǯ�B���{
J�e
��f�<%�$8�Sl�&����_A�(����C᮱������q$Hsc̶��9<^q��Q,�ݛY�j�g ��
S�l29b����5����]��d�*�ښ�e�6K�M
�C�6���d�����D���"�o�$����.�7>]8��]�؜uѽb�Y��+p8�N'WŇ�O�@��?)ab:�j-vE��k˵8/�&��F�&+3�.��e�1��Y�J�	�&�^[����#k��ɂ���[��aV�d��[j�4.Ic�~�ƫ���&L]hr]h����ܛ��]�&�AG��pvR�6c,�8?�<Cq�	��βg�S����|?�(3�³��aQz�� FG�-S&$��c���b����h�P��.SCz�0�!���?8[�UM;��'3� G���$�J,����/��*�/�fS�qyy��_P�X�ݮ�v�l�w����U��D�X;�5��k�l N��ar��¢�+�:�9[��`�U�fÏ����U�Qqh�zQ�{=�ƽN�x�����D%��}J���n���S�C�j`�6&z���q�;Cw�!j�˛P<��ĉ�"*��ʏ��ϯ�}^�2�OIN�{�n��h�k�6�{t%�*z[����-�ʻ�r�N�ΐ�1�;�܁y��_�_W�f��G7�"���3��<D@)sX��4�^h4��Tq4[��]^�rm!j