��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�&@xAMhֈ���z�	D�ɴ�$����/{҄hx�3�C�[�a8y��x�y��#sA�+q�d��"��W�~`I��|�t`�Eu{1_�v�1�8p��c�}O[���	"N͖@�؅ʬ�̇l�:u�c�u�6=<d��[x�f��s��BX��Fj�2�4&�KA��.���h�<5U�f���2F�ˇJ/_'���Z�Q3�H�)ӃC�0�����K�$���=H�\x2.�f�a��w�8+�\}�`O�r�~���j�����~](�907���.�"�mlt���+�����h�S�~�~q�_�{Ew��ή5}E9+tr�S\{_�%7����n�H��SYr���-����覙���M���L�A&��*/�����PG�.�U�P��;�G�ש;��\>Y���k��H��8�����r��ѼZ��A@x��)cb=o�m�`Yʱj;�D����;�
�B�� �������0l.�/Vl8ƙq l�\�)��#Q����޳C>|��N�g���5��hD0�96�������Ory�G������YX�LS;�6���S*��B$�K(@��toӥ 4�ϭ�!�m�>�<ҖQ0�q��\Ȕ�����#p?K硎k6���>�A���f�����ezɿ����ܘ�!�%��(^�!�]i	���CT�����4����}��.�f��UA�Fέ�=�� -�`p���ٵ1��r0�Xj�u��@lR(��Z~��H2��#�� �#g���
r�&���N떾 ՉJ2\_��Zg�BM�!rk���k�e�@�];�P����B���ā{���v�C�v���gQMȥ��\�C/�|������$8���h�gpd�Rv�Zy:sz��xp�W����|��\�'JH�y����"�8s�}���y5�@T����.�F\ �ۚ�`ӳ�D��o7�k����!
0�B�+.Ȩd��K�پ�Hx*�H�Qr7��~���𡎄T�h�f9Ѩ���8]�O����9mU�؉��5�����ۖ�������ayE���6j7N>B�D����3}hP8���4A@�7=�z,��ԂU	�d֡���g���6���i$WDpۺg�Ư�� �v[�ҁ���:�ɠ��N�v>��2z�(>��{q�{�n�,��?ϸ�>,�"o�=�~*�F�j!A�J���]��caX�ٷ�� G�b	�[1oo��!��g���H�j(gna�N���M�\�ěyuczI��t!3�ĜIb�-���sh��[���%�������+-B���0fCZu���jY�!&���^r�!��L�5v���ԇ�|7�2��
�M��@� t}���]�5\�Ol�od�➈Gà?ِ��g�	^Tx�Ŕ�q��)�6o�nb�Sb+�K������y����$�=}*�?��]��2M��3��ߕ닽��U0�Y�!���>(u��f�\����#=b��,��#�Q�B�9�����[�_W���@��m[m���.?�Y���ɰ_��ʎy�¤�z �N'��t=�&��(a������nC��褨���ckh�@� �
�$)��<��֖��[a��n�SR��+����e���j�%Ш�����	�[r}�f���v�����`�6����w�YKS3AhJI�PB�(_����o8���'����I˨!6��$d�^�C=�Y0߃+��c�|���va�.��n�&�+.����pF���%���*Q�d���ʔT_Xj��5��L�N�2��2�r�j�kY���0�������8����&����u�r0�y��3�O�)u�=�`���1r�!wqimA:r	��������ނ��?��>���b{;6D�y{�vKٴ^`I��SA�Y�-C_�}$b4�L��nߑy�oOV�Q3J�f���;{�9��X��h�)�z���ۈ ���3�IVլ�9�j���Q�4�f'�����u�X�bk$���7�gK2��,�#4��v��Vx��64Q�0��8,��e����YIvC��\e�����"�d�!�I��5.��~�O���9����Ri&`���R�^���V�:]�T��︬,E��%������CH�ؒ>�h��T�.���s�tc2�+��	�spz�Y)
2C�����6�.�%���L��
AD~���O�Z�؄I�x޳h A�8����n���/����k�Y&���������H��� Z�Pzyԅ(<X4e�މ�N�TH6�S El��ޢZF��EU��d������e.l�6��H8k2	����<�zX}h�2�1���5L�1_^͕���j=,١�\&�Y��nEc�=C1pֱ��}|����hA� ��H駿,5y��ҙEճ7����2ܗ+|)/��%�T~+�U��>����%jy���ڸ��HLd"T�����wmKC����	��2�Р���pSd���Q�����:�V(0��Kڹ��ێ����EZ�*��"���K�@��vF�r��vT��=gSn���&ʣ>��5 dm���L�V+U<'xgP��`e�d8�*
��������5[�o��q�b��N�,�0��J�(н�1�V����4!��$�n��a2~A�����vӶ&�:Ē�S�^ �����>��M�)�OM�����S�#�ɃQ���
��Т�w� ��O���ryC���K\�J��,��,�>D�Q��~G��ӚF4<iϹH`q=j�:�1Da�&��:�����i)(�E��.�<-��1q�#4f[�`;�� ��Dt�+ouخsל�/�#5�* ����]���;�ӟ�0=�{
�[��f%�����J�B��$zs_�������_�C7��}뛙��r����lוScN�d��4	�_V#$�M�!�l/�0i�^�����u1Ŗ�=���}��Do���<�1�(�p+zw,�E���-��>�o՝Px^�գ륑$I���{m���DO�Da&��c��i����p%�>;���ք' `´���%���pP���;�*Ef��h������Cz�w�\"�=�`�0א�m�u�F�X��c4��s�������ʇ�|K�h_H�ʇ����>w��nA���e�(����H����8�e��}���.����'��m����,j�S �6�#�P�zƇ�-m
�-"�Z�r\@�E�ɖVY��Z�G�T�5��F�LV���]4�ݐ���!��:K'��$�ƿ��P�l2��%�ֈ�-'�@U��P�)؜����*K9<�6���:�|l&��Ja����#S�W��Љ	�:�P��6 O#��^Jis�~�b�v���x�Ȗ)哒�=�u�F�b����������.$,|�ƅ�庇K2�QsOP���lc�ʷ��_���-��Ĺ������%�~�S�n�d�˛^I�up��J�LC:L��>�F��-�u���@��|q¦-�c��x=����f�{q#.��9K�5�*[!�<;�@ĥ)+3'TC���Ckw
~����N���T�F���5Ƀ ��X�p5�.a�]�[��X��^�C�A���E~���2ڰ��ﺪ����fq��Rh'b�[q�G���Q9�8u����JW|d�'�~�mOԃ�=����n������6��� ƣ��8����K�W[-�����]Q?����:&���y�Q��#C+����۹~m���x6~	�t�S�����cԭ	�&���%訌3�ؓش�:m���g�f'���f$պ�iu&ypa9D1�^'V�+���zYXV.�}�/(�)���b�|���J#����]�=#��
$bK�Q�����Q'���l3Hrb���d�#p�EH�ɈVY=E����(c� ى����tMj��+6#aY}0g��&��cO�WJˢx��#V=�]�|�(���S�w��oW&�����.Z�������T��$�	�\�UT�aPl�V��y�
���l�$�#پc���_a=/��L�n�p|aO��)���A$�nr���;��
�mj���$2�Wc� �JX�<��/�s�mG����i�k?!�k��J*��ܚ�R�v+�a�A#z�4��®-�:7RcJV�E�ἀ�ғ9����P����#��F��	n�0����+�fA��Vik�^��pN����{�x��hx�c�:�����m�l�G!�Aȏ20R�!��pI���r�3"��������uj�(m�ߦ�a�׎=��l(?U���x�W���F	��ՑWa��Υ�N|�������c�q�1[�����ҙ�B�I��$��|�۾Q��ۋ�҄�g$L p��c�W�G�V��|M]��v�i���o��ݎ��҆���Uފ�U��K,oi7�=�m5\L!L��~���1�(��5B����Xڈ��keMݍ�,�$hK���9��0NG���[�EM��5����I�G������5�6c~��S@�׽FG�g�d�'XH���"���*t렩'��颧��<�a@'��T��[Răբ̖K�~��r��8�:C;ƶ�`��Yv>O�{�_���"�k�s͛��J�P��R�e���$��a�M)o�"[�֭�S$O��͗P �0���6Yb��_�jD�&��Q,O٘��_Xf7��
m�����n�F��C�:�O�٪�!-
�ӋB;�}3{y���`�ۿW��O�=��Ua@��U�Gݭ�p�х�әD%��F�L���k��G �����5x��`ú]AhGq����u��A7�/��OK���߾���@2'��)��6��L��ߎ!�u�o�DE
^ϔEO��g|�XZ&���0�4B��uh`;��-b�p�U~[��kп���C�eXm>�����HT_e�t>���<�t� #+$Q�5D�0��V{l��j�y�Q0}��%����=��г�	��<v�7J�*'d���a���ܐ���T���)q��� D�@:G��*�n��M2I���H7�V>q��gJ)W�
V�`�I���1�Nv�Q��/+��<�_��a�R�:ۧ�Fd�}$�OX]ԃJJ�4C��em��e?�R����S�\ViK���ɫ�����ő���C_F���(�e���m�2'RV;m8ǃl�1`��1Iw�� �g��i7$H�a�H��ܼ�cT�	��Q����T���N��$�F�lY�3�뮢�AI�!��|����b���nj߬���Z*K���`��3�H�[pw<�AU�-M�e����pV:�� |Q:�ur�~>-.�33�R�e���ײ�ENհV��fbrd�׊����E����蝭��:��hʆ�lc�rl~��Dsk�8`����������?xv��LLS`�<\O �6�g���^ܢoh4��Y����H���w���>��c��7��e�N�I��Y�s�*Fr3��ېVl]�*�}��_���7EA�����^�׋}�)�1Uo{t���c�o���-��]V�֯��p��-�p���L���ǿ|�p�	Di:Hm�g�#_�y��J~��[S��P���t+�ҫ�A�sUo��T2��0�'�+��Q�e�����<�����,vtn�Y�#���0.rH�,����f�g;���bTV��O!"���HY}�/
E)�1@I�/��m;3��6T�G��h��y4\5G���k詃���ĸ�]e�27�����Pp��P�P��?��c�dD�d���= @�%/L1�{���^�sKm�X�9�w�J���d\{9�'g�z���fH�*�X\k�?�g��ilS�i����B��?�k_N�����h��!���s��-|�?.����c��}n�.���4�����}�z�:c��G��'`����5ō{m杮�.���!�,�2�g��.��#����kƮ w5��Ӳ]Fq��(�N:�iG oG�Ki�#����(��1X���E��v��I�9JTE��A876}�3��/= 4�Z�AnHb�F}�6�� ��ˑ0V�<��U҄6�B�-�>,�'��%r��ID̫9�zH����X�'>%\N#�������Qf��	����1.�q�ȎYp-�|�<�6�nC�W�����2�-_l�h�R�l���T �x��L���v�Λ!�Wnԫ�!�'������jHa����|�<�����K��W��5�{%h�tox�ݑ���G�68<*�T���˽��{��_!|��5S��?<#&����Rc���a�h1%�]�V�7����;M�]� �K#X	EN[6�F�|�g�|����-J�$;��� e(#Ie�	��D�p]�q{
�4)�Bb�۰������Yx�.,'ϯ�bVz��8��{����=�T��N�R�Ou��!�,9�:0���B�����࠶ B���@�+�;��$�& _�C	��������He)��5Cje�����f�^/�|���e5pt�=�@��}ι�8���ڛ>�)���>7������Z��ewΟjד�Mp��ڸ}Tu�%U�R�o��*UyB9;�d3�t�*�z��\뭙P'�:>Zv�t8Tg}G��2ퟮ4�b:����H�¨�3���,2w#�?h�<��Dw��˻�1M�FXȎh��F
7^��n�?Ɋ��s �g�����9_)�qm�5�8g���	@���[�eoޔ�<,f�;R�"�U��2a��n��#��j��Rk�TOj�	���Y��m7|t�o����@���\� ��wX��ev���r��Hrmx_�:��E��M&M!����pF m�g�N_~(Hl�-�+�	Ml��/�O�FYϙ.��}X��	_z��rP�D���&c���ξ���e���t�?0q3g� e�X<KM9�-BD��i!����[�*�nX�u4����rb���d�B@�ہ4�^tO�}�X��Oܝt�ݞ�D>��fC���k���|D�;P�����z�mFDX�`�g)��y���i��z���A]�����Շ�{qǫ���NG_�lrD�Q�KP(�A�����@t��y�6K�Z�s7�ױ!�
2��N�4��v�H�pk�1! �nj5nJ��{���e��v��bKQ���"�o!�4�>��"�\���/�ھ�m�f<�rE�巩T�{S��X���	��V��� +	]QX|\����jeC[�A��[��P��*ğ����|�7BDݔ���x�#2�o�h|�����ᙸ�T[JF(�w�ɥc��.���0��s���@������������J5�]����  �k�x��^E����'(��J��p]11F�����z���H�L;@le�� �\�FN$M��m���/"��ֲve�*�_n;�˨��<�ԋI#�V1�7d���b��^�]>��9E0Ho<�c�$�[��CE�2�o�. ��}����2�~C\����l�[^�f�����������Mz�GE�c���|q�c?�k_8K�-{��hb`�Dz,���߾b�����_��:����_������.:ib�ƥ��'O~mSU��Kn ��h��Z�?����.]=v�L�,[�������El� |��:��p/�FXg��l�S'��mR��;p���7�}�W(��L�>f��Y�6��@n�@��Ks�1�G��1�#�q�qh�29����K� 4�$U0� �B�� ���e���W%��p�~x�1��X����m������{?V���Q�%j�h���R"��<�b�n���7b�)D���m*u��%~��4��,�QY��9��d��^?5E�[M����j��ye6r0/��SK?���{ǥ

�w���#��,����������f>���H)����X� c�O�����#8�qs�w`f~�V��q$ɣ������C �|�ý<�������y[B �<��a (����cVF����fG�V\�Uᯖym�a	�~S�]iL�����,��ӛokZu�f����{WQ_6L��[d�E�]YD]Q���鑑��@�1�:˾
 �{�C1K�M�'ߪ�T��v�"u�<�l��]9+�4���
�mk�"���������n3DJ����Cl���!Q���vd�]g HSn��V��׆~�jk��Hs+��66L$�k@LGb�i��������_�Gd���4M�4�M�ϖצ/������2Ƨ~,E����E��^?��](j��g-f�'<ϳ�4�)1d���h@���5,9���9�Xi�^@���邊#:_z<h��{S���jBGM�o;ѷ��}|}m��C�=Ҙ����Ƚ�C������cq^��
^�ґ�Ĉ�� 
�L�d+�ШIebSʆ���>T��,��%���*�D�+}���p=e�xCO�7��'Ǵ�v�����"�P�3sD?:��GJo��?ixvꅆ )�|�}j̀����)O�io'�nL%�V,�M������:U�㹛uʹb�#"z��Z���+�pФŻC���������9Ҽ*�%�妆T$�F}�$Nh���N%�s�((h#��L��L�]-�	`R;�dY0�np>a�jc�L�lt�ɝ9�hK�+��B���١�r�x&�h�����s�h���g�r�q�624��a!��#h ��cÛ14�*-�@�k�=RJ��V�s��U���p��f��BeG3��#��h���"t��^i�y��*����Z�uv��=�gG�����b���!U���tĽ�f�6���.����[�:��p�R��,�昚��ZTU0,
�ȮD���be��ހ�k.W���$B��v7<$o��Q�)Fg�_�q
�b��h�ڔe|��M'0�|��c"�u��q�_�hLm�Li�r�#�8�q�TH��7��Gq���<<��!x�9�T�D�afz8�uu1$�PN��`�@˂T�3��U�=��p�s��rg/MФ��^]����{�/�>3�.f���t���ަV����_VIa�y�h�x��)4g;�_%�ܭj<	s"_q��~H�A>Ӎ	��O:�WL�6��s/>�)�O; �pj�՟϶�N[��2�>i�H��fMh�u�xy��M���u-l�Y��0!�P���8J�Ⱥ�J��z��P�"���+4�q�ۇ�w/�g�<�eA
	a�ǙN�I��Uo��!���aʤW�iЈ�6G}��h���<u�����H�����cTUZ�����������Lș����mQ}b�땒���X���#y]���}�2��#���˥�ˀ
1�k�qXAܷA�|[�����P��	n*l�6�P� ֽ�	�#��Ƌ�ԙWSӎy>����|��GB�+h�T1 *�f�y�r�ox�L+>x��	������9ʍY����ث?`!Gcsm+w>�%�k�&���򻛚@���yVP?�V���go3* �;rOB�ې�����P�0�6��r"�Q-��%I���bBZ�- o��DCj����aa	�� �d ���Y���<���<�T��ج�Ƴڨ*ǿ̬s�#�Q��1ٷ��Ȣ�n(�������$a��Z���'lʢ=m��xc	��t��.#�^����,,-�&��O��I�5�Z���*�r�Q����on��#~�|����
�Q�D���k���o�j���ɲ���3y�o4����\�Nm�`?� ?��9}eyjU�&�XҲڣ���WT��îʥ;`F��4m�����E��k)H��Q;���LP��-��kd�C|���8�g�BR⺈�H��{��(��L�}A�.�T��{
�VvK�E'�"��H����ptŁ�p�u}w��=�1~����m��F�ʒ��n��7�I^��h�P{�Jy\��k�mIMk���2��kԮ4
#<!vR�B��ـVO�ѣ�a+B���
������kk�D�`$����ŃYL$}Q/���}��De�����$Vd�-�xD���=o��cFʹ�u���~�ϮX׭W$������
0���gc}�f?8�-|�v��h�'jiyg ���zn���qT/mwS�����=p��W�<$8���C�T�ܯØ�3۴��dP�[}�Sf�ý1��8V��S�d�3vBկ �H4
�L�s�+^�R�6���[� @�g�>T���f��g@�<s�U���E�Yh��O�٩
!�k"ŌB[���_����rb�[ȶ%̍O�<n�E�-���ٜ|g(��m�>�G����B���ؐ`��'�k��gH=���^�Әꪎ"�,Vؙ�c*[�[ƿ�ޘ��et�p��(���+�Ix�'���!~9|?`�"W���Pn/�kA���;��v^y����G�R������%>2������LM�;�ƺ��Ys��",!4�5���a�s6���/��ﶩ�x�B���]��_#���opx���%#��w� cm4!:�{�4���&>�a���-U!��X����O9���2��t�d[2%k�|��\^�
�	�N�^n�{�_Ѓ�@>0��R�jDy�4U�&1 �d%��D���ÛVj=i�X3x�D�MM�'1�wԵ���e�oQV�66>b�L�<7)�iл�>��V�}S�ї���Fn�B ������*ݾ�?�!��W��6�W��KS�op��!�K��6'�C�P���r�Ƀ�>�*sCy�A�)Ɏ���������u*����1����"���+��m)m-T�\:���V�7��qP�z�s��n�I�xH�OQ�Ϧ�Q�
� �#�G��S#� ��7��b��y�?��J,A-����N������,�m��7����A|ߝg�=rY|GǴK�	P�&��5��bw-h��?;�����g͔&��OJEd�n�X�ay���'ǘgH�2�`����+u>���}R�(�ov5���?xJ��OT[,)�b�LK뛢���F������7^�ߡ��o-b�4W��ӭ���>|�7��|&�aCc�IϬzƼc��H��2�n�o�q�֔��͙O�uWzK0�o�]�`{����(N�Zt
��ah�Q� �VP-/�{��{�W����@FM拪�� s�#E	�u ,@���W�w�ӨG::� )֐��H�f�ų�y����JY�f�[�J����(_�2�-�͂<h�irs��s���T,��{�QcpM��'D-�Q[��^%��9W���Խ�SJ�� ��Q���Ʋ�ϔ��*g:��4J�{`�7]U@[��.���U���ՌI7��\<΅E��Ɂ�XZ&���Nt�����r%m�x˙tĲnUd�&KQ��>�{O^�f��?G�\rf+���@�a��t1]Y�{7t@'_;,�zwg�60q��!��/5�����F�t&'���M�Ja>�&�-�(�����0�P5�!�P.��/#��Wʊ�ǧC��B�p	�Wȧ�����/�#�ܑ��|J�f�JT�4�я�q.���D�<�q���I^�K�.�zN�5�WքGu�M������xC�i�~��W�K��ى�iE�J��z�[���p�9��,�4c8�x��wfda�`m�xNݖ1���+eD�\3�T^I�e���03?o�m��iQ/��Q�Tu�΀l��t��~��<v���n0��֐�tֽ��&ຢl�m>^'�2��:z�\53H��к�I���]8�P�6��� B �E���R5t�5A�J9ڗU��V�';w�C8�����Q��$��}��J*1,W%�_�W]S]��B�	�ɗ]�wԵ{E}Q_(l;A�kMwS��>�����?�訙V�13���Z����� ~"��B�����-|����W���w��0�*��H�i��L)�����*Q�H^щ(G��;�С��U�#�hT�Cr��eޚ����������ȏ��.4���&�s�t�1��$�p?fd�Y*p�H��<�:�F�,��߭Gd?idf�~NR{B-m6!�-g����w��C&�q5�͟��Yz���c�w�A��in��� a�E�~����횳��Z���gE�|���؟���j}���ǉ��?�_p�($7�rHJ��>�~a�S۟�%�t�)Ħ获`@��p����*��c�?ؑ�����<�%Ho.9q�|q[���ᶄ(�R���侧�7�􂅢z���|���p�\N�x{IT�ǂ��_� I��8�k�<�?���s�����+�o��\�A޳hBm@�?��:��<y�����D�"�v��w�B��c��:KRH����]"��=�4�s�7�vx���'B�<�c�E��x�	i���9y��k����]�IZ]�� L��F���g��l\��V��F "���X�#d�2ǻe%v���5�Ƥa���x?���y8����u))
��#���GO	n�~lXU���*}V�3i���
Kz|�.�� ,wr��=A�R*�
D=.�m�R�8��t~c�.���^mg��	��� �	|:�������5���:e��]~ĺ�L&:�ڟ01�y�"�ge�o�U��{��7�nV��uv����#�`0��H�-C�ϛ�m �,+=�*��G��ލ��i�-IϬ`6B~��h�І���B�w��&�S��a��PѨ-���"����P%�R�I:�1��;w���U��>(��:lֽ�_\��~jҬ�a�P�n')�E��m���9�ѧ6_�a�B��x�"Y��Z��:�~���0K`�E���R�:��N�@؞[�� �K�P��aԍo�S��|7�X�;dݏ�t��n�Ь�X58^L��6ig��ĭ?2G������%�7p0u0���jZ4d 
#�%V2�87�-����܌��z	�G78Q_��#�M:���'��z�K��}�<��%�l�{�i�L+^������ �R��wj�q�fn�<�9{c+�~ofPm%k��1�U-�����|���A篱4c�Gv ��H$�G�< Qo���k�)���V�~���H�1��a�Kp���*��r�?	�hr�[2�*%[b!������K���� ?1����F/���5^�/��`!��D�Ϊ��yL�D��m�-��?%�G���5;�ρw���[�;���>/V������G��wXv�V��l�	�[_�\_W@Wι������T��� v	+��}� ƚ5oq�iO1����QS#���y�4���]�#(O:@gK5N�ଘ}���aΐ�����0�:��_��M�\�5U�S�)�$�#	i�]�J)��)|E������<�'ݖȲ�}���ՙ� h���%4�D�U
.�SgcQ	�ټR�P6}*�x���ȗq�T��A�V
by�+|@n�*�%�8,�b5�HQTJL=A��"�COS��Q},D�t��9�|� r��'/ß"f�)��2�ԹHǔw=�F�<ׅ��j����]�M�kI����ƕx��P���7 �˨Kdy1 	��\2��p����xC�4�Q΢VɆ�؉6 �#J�T�F,�2����0����U�.֝��4�]O��?C���8�Ó���
_����8*#��\���)� �ڤii�u��7R����q}�Ŀ��]�dq�ZxgMG�~��h���G�G�����W�����m�EP�'ߞ� ����'���(��ͨ�Q�Nbғ�XE7*K�7z
X?�Z�=&&=��0ͦ��N�Zr���/,>ဉ��rn��au���[���N |��3�n0���2"�2`�§?K�9�?�hF��#ތG����U������P�2CiG��*�4�D�ھ���X�e�3�� �zb��y�h�o4A�JT֚^Y��I��@�_b����V��0��� �O5bKV�M��]��zI^0w��� �� ���z8��(��>jﺐŎ8|���=���=�D^G��	3��pQ��b��N���� �nAJ���F��/�$=�s�:��) ��� H�� lv��*RC#A��]M-n�	�tR|�)���nr��!�s�G^������G0�҇ ��� ���h���!u<�/eȳ�>~w(�8�r�3�T��E(a���9 a��t���	�yr���b3���ĨdM��,�ߤ"�[��:�_��^n�!櫝 I$FIek�H��K�r1�9r.V4���.e��,8#�&�%����!��GBi�'�:m�ы���`L��o��˯p�_��ILB+:-4<wi�M�^r�M@����(Qq.2'�c�>y �8h�{
& h�_[��/Ce��K��!����7�֬�xp��:���'�ۊ?�2��zu�3n�jhk�$\��d�3����v~���ZU��B~N���j����*�F c��Ģ�h�ҷ����$�_� ��*#F���tKy��ѯ��ܤ-�p�#��Hsد r�6ݛs��'��'�����Ì�d�fOD�c�E�J��7R��V�)����л�X�<���rֆì55L�'������~��)zT}4"K\�@ 3��k3�u�T�������T|�~����	���w@`�b�b�>��hQLau�Ĵ� ��( ���9t$o��=h:j�~�Zl��l�Fܘ���󞹉-����J��Pn��=;f[&�����hr����+��Y����uxz��d�Z)7�f�����B\�Op�s�ꋏ�"I�+$�{Cjb��M��c������� [�1���;�L�ީ��\p�c�ԗ>HMk��0 ��w������wo���pT������4�k�˲��o@;_��N��K#E�X��Et������d3X�p+�:5��&AEx?�����*r�j�xE{�fc7�U�UJ����!nj���orI�����h��ݻ̐������lۮ�{�y���>=���&w�tg�Ģ��=���Q%��2�L�PD6>�fW�@�/;q����N��dZ�M��鎌�1gZ��b׌��&��j�'�'���99I��7V�@��Wȼ�Aql�#{t�����O���-?|eB��RMu�¹S9"��&g�R���n���%F�n��d�[[t�a8$]q��V��1�����<��Ϻ�d�I�ꖁC��4r��w����o�8U		ˢDI]Pj!��u+o�ĐE\�
P�l�	���8�{�5tz,*!��'@��'6��lP>
*�	�03h����:���	uas{��Y��S�c"\3�"m�s�~4�ߊ��Y6��$U���PG��͕L!U��1A�S>|�)
�"LS�Fm|rj�1�S�`��Q�}�5��ca�ˌ�7��s_��)�%�YHWI��z�S�ƛ!i���EI�c0��Y�~R�L���7n�u��~�|�h2s7�+3kX�� /PsR��ZF�++bk��Je�s}��T��"�V��8���� �:ͨ���hq��Q�<����?{]\Q���ay�3u|��F,dE�"�D���g���$6�a�Ӭ�6�Y�f+](�^6��*Ep-�l�:��#?�����ӛ��טQ�d���І��?��?N�VM@�(�-^�]�������[4��&�l��q��5L�$��Q�1l��9�c��RN,����U��2�|��=���<�4ڜ1���Eͼ@����AH�A9�b��w�_��3X����I�6���fG���X3G^�v�lQ3�Db��
y��h<�Dɮ_1?��#��K��������Ncɗ4��,��c)Nr�5�)0ߙ�w���ٍ��,Q�ߺ�w�_C�2X8wlW+?�:�
#�t�͍elc�����*��Q&�^�/jZ�w8����[�R@I{y��L�'�L��B���ȉ�d�ӛ9��7 J�����T��V���l��7�VD�	�G櫆P���jN�� \���NP�i�&�:�N���.���lpԫq��'���^��ү��ӳ|ԡu6np#�j��1��/9�!l��۸֣�dRD�UNY���������۟&�仌�F�0�J<����(�)���Ɨ�_A�7�*ŝ~5(����>Hh��Y�>��s�b6G`�q�콙Ȋ#4-���)�gѩC��$�ߒ�c�+ܦ��1�0�����I
��^w��r���N>�:1�b،��"�qY���$���q})�<�@�1���1�?�@]_`a&�N��gQF�}�K0;�gy�X�'�ߖ���8��4���
�����˻X� �ؚf�x�[�݋c@\��/�z<����{��<�Sf�Q�������ߍ�Ǐ�eZ�H�L� Aq
���g�y���{F��$&� �쬛D��-�*��
LF"(U���S"J��o|I�M�gV���t�i_��N+��߼C�OK\#����3j_�����XO���P�?��<���b��j���8�_����.j��K�e���,��x�n֋H	���t�O'Yƹ�w9������YU<|d�O�(�N����Qi�r��p�����M�rj] ��"�-�=cq���d����3��ؑ�k3�� _�,%�R�/����oM�cQ�!�����*�N��ϭ�����B(7[{�Yԁ��X������L[����}ѱ��x����Gy�o���0kz�(
U����v:	m���ǉ�a����8樝S�����!fˆE��E��=	�k84���Fgk��
:����oF�8�a�Z�}um���N�lh�n���]χ�������cQ|H����@.ͣ�H\r�Y�m�mj�-�n�tZ	<t�9*JB*3nP���?Y���pק6ab��>�ƅHI��D}<�
����w�g%Hd���e���<���.I�~���$���������h*������(��Bp��\��7�Y�\-R�.~�:�J3�<���KZң�zP>�pa�KK[�dO�d�r����z��o�L"�j�m@Z������n�{C�3^;�}�[�z!�һ�!O�A�!0�-I��_UJ���˦>�f��:�u�X~��}7Kk��ٖ!z�'F o-�4��0��^*�pf�A�²����&��3�z�%�o��K������>�Pᕘ��b�X�4����8���wn ��Ji�p�nm���6~���Ù���nfM�|��SYR�i
����+����d]O�Nݝ�{[��z�����
x=����-t�!�Q�Y\����II�8�,���}O�����yA���j����apG�wC���ҝ�y�dIw�;f�A�yG�+5Q�����g�bW|�y'T��a��
�Ar�"]�;�g�3�� #��U?7�ō܏+>!�P�t�]2v��˜p&Y�+I��&�C��OH��6�����K�Z{����VC�mw���-���ᕅI��\�	��'hu��$�H_�z��ž���4\}����7� ex�RVwhB��\R<��F���L'�S�`��_��g�XːX�9�G{8gG��2~�A��ӿ���}�G-3�l^g���QB�Z�)�b��3����p'ΐZ�ҟB�L���A�=ӎg�9o���SHY(���M�r,�ͦ����z�MS�C� �o�K� ���a^,�C�>��alD)\�_XUf���y�6G�z��׀;2��y���W#*�4�6��ݲ�
���5z����!�(3hi�#�|r�:\��H�)^�*RѨ���L�B�|U�a�HC�@�KHwoz�3��<���q��<�]�=�8�=������qX�I�6��S���b#7�
nfޟ�|?�~Џ��Z�8oYK��!�� ��ܩ�#�'�e��%"�}k��������7g��5c����S��I�3e�����@�Fw-B��K�����BH.���'��W"�>���^����Ǻ{ <��H�2 �H�*�4��[=�Y-�k�w��%'��%h�|��q��4x��E�|:��2+���Ʈ���^��n�m�V��6AO43?Yc~%ٻ-�旹a�W �w1H;tԩ��`�1#6�k�%S#QīN� /�'�h;ⵖ��gwm!���wPO $n6��w9��O}�䛿�LT:q���cÐ&o��9�s71�T��wb&��}�������uĖ|~����WY$�+�'˲F!|��}���c��ԫ�6� �(R� ��YL��v{�D���ב�WV4o������%{���
�U������:0k��% I�^����a!0����Z.ӛ\j
��SΎ_�-Ͼ����iߟ��o9S�
�0{��ŭ���@�H��O���[��@!����B�Zv�z�zA�|��Q8b&	�� 8?�v�9˪��p/�-���l�L?Byn�ri�#�L�*.�P��#T�&���q�I�Z-C<��UPZ�Ê�|�QDr�&˥-���ׁ�m�O��c�Ȍ>�d��;�s�*��kT"��B�P'��-E(��2�ɕ���A �����猕������"L��#g���?'iL[��<�h����yO�=�B~���\�
8�Z�^�9\"s����S��� gt䊨�x�ݖtpbFe�O�A^�;p4ڡ@�$���t�,�1p�������p,�i���1w�v�JF��*Y�`θH�� ӕl	 봪����¾���
��8S���~�����!z�|wf�جD��*�x���M.a@�6B���=+�`"R5���mCjJ���	z[��`�:���>���|�#��Դ�=0���b�ˮ_I��W,�΃��JB�1��h��B�w��S�OE[뉶�?l�u,=P�>�ó3+�4E�t[!�/���Ϥ�9Y�t�G��YS��'4�H����jbO�g���6�X��S��<�P��Z��/����\�Ɍ{��=)!��5	�"���CU!f*�izHɟW�呺�8}a�ǋd��!�9SiƲ��Fj:��9;/F6೥�Oa��ʗ�� � ������� �����j��J����.<m&Y�-u�u�Ĵ���fl����[@'�Y�Z�fO��Rpt���TvB���Zy[[��z��n��_��E)Jc���� [�v����%�'%��d�P҆��XΝ��tf�Tt����|�?�BT�@��TE���D đ�X��h��@���׋ܻ��_�F�_8���J!�d#�az�>�įgLq*hL�3B��9���=V���Ԝ�3X��ք�>z���P��OzQ ��c�^P�88t�:��F�z��L���al$C���GD�:i����[m֫p-�����q�x�d��%��>���%���GYc�l���F�J�KY��d%��kpfTՋ�z)��5�<L9�7� X���ʢ�Љz����m�I��y�k/ǴH�Bc�G>�G(���r��7�廘�^�~�e���D�`��k�� 9�h?�<@��������l���$W�3�Z�ʵc�+k0��@������$>��G��qn�~��f�\�$��}��&KϚ��rޟ�.�t�_�B�k�^��T�.�p+{�&���̠����?D<˔�梁��_����H���k�H� ;}1�4��Tw�����YP�E�\�g��s6>'�B��0!��������懚v�&+s�L��|?n�T_xɎ)i������4�_��(ƈA���,�����P���t����_�4�~�8�.`��%�S?к�ÿ5�6�3�����m�<)xГ%�ve*[Tu-5��r�����N�g[�;�іW!�u^WU���C8�|�*z�d�)�uy�a����N�X�6@x$ ��P��T.dڧ��E9��֦� w{T��j�Uߧ�OF�py���ne���̩�\�D��r����v��6��{���z@L�� �`��-�H����
q��fɅW[W�1<ID�p�"s��t�a[Rt��Ѫˀݾ[l4$÷se?|�#�s�3-�܋vcك��2�6�pFЛj�Q���x	/O>p,��Z�]��2�a�)�#������h�}-�XI�bP�l\m~)s(p���U���@ڷ߶��x�0���I��@l�QDeF05lf�¶������_+o�^86��Cڣ���Pη�=$�W.��
�Z<.�H�1�L�I��H��f�o������Jd*�8@��P���q@iE��~ I�&�Pm��..�-){����U��ϓ��>
W�� �E���4��ʴ�V�_Ʊ�e&�M��T���PBqr������G.��ubA�읟�!�`8
Q�G�Ԡ�}���bY�jI_�� E�,eB�;�����,U�6����HW¤�a��3��"a�S/V��0�hk�(�@�?�0>�m�	�>�X���ĂV}���ݾ����?8�����_Z���w?'��$�Z��JCM�,xz��G�n����T�:�y��(��H���Q�q��{?<��m��_B����G9�Aa����kԘ���z0g�h$��"�o���{<��\&��$�Au�l�J�
'���h����uo7`{1����ɏ����R-��I�==���5�ZM�3��F'�zn$f�¯��k����p�,�*D6�[��׼O`L�Y���m�Ψ�����b�zl�lAlë D���9x�<G���h�NTi�,���{�G�+�%�a�g�w��6[�C��3r���&�(i*�@,+wb:�����Í�W�G�5	��;��@���%��;�{r�V)
��n���BN#�1>�n�$�C�:�&:��3[y�������1Q���*an���C��'�<K˵;��i53J�GWG<ꓔ~�e�	��3����N���GS
;<߫�(6�o���Y�v�<��a݉��=�p���ѸZέ��00�'�$�44�����߀��g�����>C�~���]\xn���h��K�p�jHS)�/D�8l�} mQ���c��uF*
�!�y�0�}ܴ��(�УE�S?�EO)�c^`���8�u��\M$���|����z\Y��t�t�����Fg�O	G܊�k��m9�]k�v�w�PG̀ݤߎ;���Ӈ3_�ֽ���7�����8H"WG�D�oTM��O�uA����U�Dc���{S�	��QZh��.���O��e̗��Ec�`�vE�$��x���ꂤ\���0/֌b�}��*�xq)QX�����L�?;C̶�5�6��۽z�$�����A��`|�� 7��о�,%�mِM��D]B[����
S�W��u�Nw*ހ�v�j_^�q� fL��EO�hڬۮKG�5��]L�9R��(����|Ȍ��8���EEl�a�O���K#��8�ՂP���[���"