��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w���>��!S��'ho)���9�D�oit��Or�/;W֋{�_��}�
l�pl�ƃ(�Z>�(+���Kd�W'�s�@~NT�>��x�T�QhaKtO8�F��e�q=Mn��Ɋ��0��*g e���<StQ�w�����N8� �9$K�|� ��Bw0������g"}.s�
m獙@��;�Z�|NZ�L5SU�N���JZm2��c�<���Yd7D�a��W��� ��P�������B�޸�R��1YQ�������ƋPѝ�	���G���y�e�jЫ��0�~2�5��؅�?K����
W��l�a*��<�Μ���Vq�4�1��\6���
@�6�彦��C˛�x��P��+'�4��F�gf���_���& �nh��n��%Y<�;~/ 4��;��!
{�{��8k@\�J+��V�����h���/�-����f�}x�L�X�y�h�j�eH31x�o����ϲ���c����3k��m���韒�Uσ����{*?���]�T>�J��H�U0Xk���Mߥ�tA�(�E��ƽ�Y�D�S��Z4�vv�)�`��P�S1it�<���8�D��������E�O��5x��h=E��j� ;^F�m������{Sq42;K�?�RA�{�Φd�������<݉K����n�mWgH� 8CQa����7gu��t�Q�ܹ�=����h[���5ďA��3��B��R�^n�kh�G8ZyJ��5���"ã��X?9��N��fj�.@<��?\>\T�k6č�ǝ����,���`�1J[~�XS�$�vއ�4��K��x��H���1k�-x2k�Vp��\k:;S8B��|���p�V䡯0�ݟy���D��%]�KV ~�Mu�_��*=_H��-�VM�O�G��H�O+Bl>�{-�j��(�D����I�
vר����z���o����Ջ"�S�Xw]�rt ]m��_�y�4�gx�.5�U�2jK�+�g�X��yX'J�8�K�/ʽz�DD�xM����t��Qk�G�gM�Hz�q�����"���$xB�w�=���<Oޭ�ҋg`Bn��.}s��Z����	�Tb��l.3�Zr�7j����Q�m���ͯ�Y�B�ȗ˱)���QG2c�w_K��N|/^�w:�`41���m��:8�Yr(��ק�F����T��_�5;�X�:nC�����aW�vb��b��B�!�c�e���_��S��{Y�Ck���:#y�j�7��?#]����_��>{�oO�!\U^v� <r�(q,�L�z<��8r�x�1g�\rCW@�ÓӳtL�ߣ��D]��m��99O�y�zR׵�U��<0D�n�1.�VQ&Z�mub�xLo���� �-'�8Է{y�F	����8�{�V��}C��째oz��c�������x�����(��C~(cV�6�)č'��L�GQ�NFȗɞh9�X�Pf�{ .�$9�D#���)2���~�M��{X������>�]Qp蒹��o�FT�~�*�Ne�T���c�w�"J��	�9Wd�/�)9��dV��>BsX��
��HՂ�l�ͩ����")���Kiv�|�߄]� �XZ����i��Il�%�������,�������5G��5�ٌF1���`�y�[_J@To�鑱��,ϱw�ҚuXW꬈�Y�j��z-�A�����.%�Ư M&zz�<������]Y�@� �-C���ﴭ�0Q�J� }��|pq�}����6o)A�]��C�b�s�1�u;FǼ�H�Z+�����c�Y�;:-,�d��Ob�ZD[	5�֡z��~b�i�_���;�`��/~yaWEŻ���%�[��	V�4�GĨ�Cs�W��<������AH=���?��!�w9#p/g��D}���b���"+ D;6`��p;?�I��G]��M0#|Ed��錶 )���߁�a1�.��Uy���Z.�І��*.���:K(�2;C>m��
"���o�z�hnt~���1��H钾������Bh�vd���f����A.B8���0�	�8��r�lħW6�����bWs���������V�[.��a��A����)k�*v�����T��B�؀>�.�,Z�mlD.y���1M�nl ���6S��ɷ�Z��!���cS�@�(���[���~+�DH�]�9(���Dǫ�y�"h�i�/���;4u˓�7�d������_���?!��J�3��X��t"�vlaL'7l�Yc||fi �&&{�Dc� 4�Ju���kx�-*ZM1,!A��U�<�Q7Й}����6��(÷o�����?Y���Gy�G��J[��XRnVXE������ls�-*>8,̯�ö�^�*��2�FU�<��Q�"�T���	�9�':�뎁�b x�y�a��.=�-���¸����SW��ݘѲ�["*�"�3Q��xey$\�e��P�Q#' ��t@��K���Xw�4�$a�SXh{N��Ӻ�8�P�Ou̚�;c�W躱��=0���3����*I��C
�ؖZ�kRf�!�'}��W�9�"�o����.�Хi�Y��<����ϔW�'ɳA�MŴ��l��2L�n�Q0�9�oK�LȞ�������)1d���ѴWT�� xj�討uV��"<=��Q����Ԋ|X�/C�؋}�$�o�Nȍ���ӽ3�z�́��լ{pV� k��]'=&���(�Pm&��Y��{���t��GߩRt��i�b�[���F��v�%4�g9��DkH:'�3������zӨ����[Ă�J��	<��a"�C�>����)��ȋ?���T��ey�wOlx	߽1D���t�>.�q���?騈����:��Kl�&�n�|^�l�����f��\��p��IopK���jǸ]0C5�{�0О�r93]Ϯ�`�@�3˷k�̳��ČM+z	��뵫����/Å����7��;�jj���e@��]��0W`E"v�t�v�1.c*���퇪3M��Wzy��/������N����.`���O
�l�0 ������K��,��T�u��<d������`%����Ic6�⨶W���-Z�z�f�ĴW����7��B�'Vg'k ��+���7���'��y�#�/�9ĩө��2��H�m�����7o�3�7��6D�}���N=�����]�k����������g�<������BF!�6p����p�q
�q�|���}&�{�� �P�	��������|��:�;���nYu��B�~��4sF$Ç� PU�;�P��w���]��2-)h�w��d+���8��� ��j,���a��Ԥ�Z��C#w�ʞ�=g+Yc����[��$,mS�%��w��M���9e�0��0���%��A���It��fi F�h8��م�XW. )�A�w��5��E
��K�hX��H�o������-v//Jf$ 
��Zh�
{:fڇK�� -�շb[p��"D����,;�?���ʈ�?���`�.ۋC�$�
�~+Ͻ��CǮ�T�C�QJ<d	�+�bX ��6��G�e�畢ӧ e�hUE�p��V���4ᓏ�;bDGAYK�ܷ�u�Z.���4|��7�l�y�.{��[��v�,$�Ӹα�x�p�E�SʬG*�kѨ�������Ec��U��v�8�;���*]�>{���bϭ:G�<���a�t&]��쟰���`8:!�>l���.`��8n�=��X�XjT�;b��u��	>5ω����;bI��)��W=�[�D���}֊X�u]��γUb~Cz�$��%���7��BP�y�z!ď"�Lm�g�W�)0-ʑ���>Y;�Y+Ȭ�x� �a;P
���\��Y�N�'��@�29�k�D(밮�/u�dNv�p�Fz�6�����|0pr΅=�U(��U��W���ﾪ1��(���sE�E{��d.�JN?�oI�Β]��~;�ku[X.%X`��_6�ol�)��f��=��~f�����]�{yp�xЫ�ח�B�0��mA%���<��Tg�՚�z�6֜�\y)a	e%�����=��q.�A<�"��&����%/�d�6/������|�} >��7.����A�[�"xU���Dp6����7G�/*u���U�L5�\\�6#}Sc(�:��Ȩ�����7mOZX�1NDZ؅�v%7��hV��r���˸�8l�>i�T!!c����s���hL������TX:���ɤ�'8}��֒'���G�M��Gu�a�2^�G����p�)��Y�o>xu\�޶�̕yh5���]���A	����o�W��AT��������W��YW�D�զV��!D�8t�����߆ �%a���2I�����iV�T~�q:z�u������b�d�9-�`T�STC��wx3�3���&SfY0d��)Z?'\�&�/����ԅS�`G<�,% ��![ªk��)�Cr-��p:H�YKH���H9�YϾ�L�)�v��}
�t��a�X����b�zw��:������GAd�i�������:5K�Tw1�qWHx�G����4ΧU{k1�	}e��BbU�+�۠U��`Q���t}�ظ��,�r��:��-h��i
fF8��D����s�x�j�����������L�5��2�m���fs�^]Áʛ"���9���a~I��5�'��)=3��0h�܅3I���
�#o� S\�l7]���~[���~�����`	ʅ�)����5+���l%6j��~�-u�W�1	�/�7��>�:$f�+�O� �7�[�!�EF-Pc-�(�%{S��*L��O�=�;�Q%�J�G�$�BE����1$�m�}������Z~�I��}����R��?�ȃj��~��5����������r�zɅ5����4-�"1�C�"g����"��&�th��:����9�5�'�F2�f$���{ƒy�ew�u�8Z�=@�?~a:#�,)�� ��/�$�aTm��>��RR�s����H�SO�o���H1M��o�E�Ɠ���Zy�(#g�\�-RBlz�+�Q�yRR�N^�ۯb4�����(�T�sidf��H����[�E*�>�Y�%�qB���R�A~���b���1��&n��
/�f�}�_	<z5�H��d����m�lv��y�gRCc"��g���j��N=�Ȏ1�;J���-�E[2��U�E��:�qOH!\����b�d��iM�@��;��ՏLl��ំ��񏬨"R06� �*�=���� �6�рU�!�=�*�"��^Σ\�$/��/ǻA������w�[�_�8�P5���[Y'Di�\:�c6S��k�M~հ�M\�	�� ��$�ƒhX���<��	輎�Ay�c�,8Mf��
i����D:B �i�_�$���j֜�z�w�!��<���P�6�V_���)v�w��u� kLi��`�
�Etֿ㋬Gx�Gw��#�e�Q�팰�,ס�O#y���T���Ϳ� -�����pDNl��Ŋ�P~!_����3;q �Ae*��4u�c'vC�ۈ�� *����M*E�P_��5�u����+��dd�i���]CbD�X������O�^͛��7�z#v�Tؕ�',��̸�ɨ�G7�줘�E@����R4�l1���_��sp�	�-����"��%�ߢHg�`E�*����vXZ6�@S2) QQ0��t|6���lO�:Ю%��z��W����ˊ��"��_�����Ee�9�i+ݖ&C3`~n0�u0�Ĕ�?Bժ�M�s�����ee7��\���6X�؁�8;�7���5��to�q�m�>G�o�vP~KoV�w݃�+\V��[}�����]��;
׭4P��$�^��A'y��<�Jd����� d��-�UN�'�8�	�.0��ȵ��O�ff%e�@����Psl�� vJߢ�IfvD ��H�$ԡ��Xj���,!���ߦ����k+�������\�3y�O����
'x��G�L��
qe��2�Su��12�7q\ξ!/�(���@]P�DC 19�
�VI<��x�y	�!F��Ff���?�#�=P�AS����w�ǩ�j��$g2�� �܄ ��p���-�o�k�.2��_�5�K�=��?��dڒ���b@���.l��_�y?����Iw�y�ܼ���5�Ӥ��cȸ����n}>,`#�u4��sZ-��b} �d�ܴ���G������p������dέ0J��p^�C�FE��8]�ʀ����P�{�h�'�Pn��i�v�b+�����˜�Qu�A-y.�֜"Іe�)Y�����R,���!�͡@��Qư�|��xM��ֈR�M5� ;-���Uk�3bqPo�1�eb	
�Z=�{W�q�,���߼T0?�x�h��l�ɞ���
���{��]kx6���� �r�<�&��]�j���F���m�r"X� ��ߢ,t쩖y��Z��8���C=���R�j��� )䏹��y�SH�c�F60��Ab�j����a:�t�$��/�߷w�蓧��K'w�^e��ϓp���!`����0�� kV.���]{%���cdY����J�� �4�זo����*gF�kP	��C	(U�Knp�Z����I��h
v�qq��Z��T�)���f>ᔥ0aJ�@1�������#��3XO�����O
�8B��i����]YꃠR�~ٚ:�K��6�?A�����B�z��0Z��~fTXr�࠮��n���ϽBds�1�����C�s]A�!��[C�kxl�� �t�@S$_���0��_,.������*&H��z%���񌋺�|�#�3gG5�"��mK��T6^u�к�D����1D���~���0���i*��A��Z����՝�3Ld"���ǆ��H��/�d�~"o��w�naWh5%�\X�w�~?��B�C`�q��uix��K�F��β{��џ�8{	̯mJ�QD�?=L�+��e�?�/������c��uYp�<*�lu9�Tj�.ȶ���F��<�P�0����cgc�#�k���E<7e�*-��J���]�����\��ݱ Ӆ���~~ϚO7#�{�����^pE�o��­Ed���W A����e�]j��� �,�/Wc���,=8:mrg�����O�+	��PPJB;���&E�����t��fǔ���2Y$x��k�a�u�,���ɒH�L�h��D�q����.�n.���
�	��C�x�s�T��Ӳ͐Jns�_�ƇAp�t9����f?�4��Ŕ]B_�6���ʯ7�)�r�긃k� A,�0i�h���_3`9�[���q�\�e4ocP������]�!U 'K�ϰ���]?؊?U]� �������;p|�\�[��8V��'@�\?}O�b����o,�ω����70�r
lA�_��x�_F�i��+��:�����:�G��t� };��Cu�f�J �cl!r��js7�:���kX�s
�H�����uzn�ê�C�ݣ�3�ػQHٗ��<��oI��W��<���B����nN-S��`cz�]��k��|s)1*+3���<�jp:1� S:-�/��[��L��\R}�L.ޕ���}
rG����v��)�����·9_UC���N�ypo}�����ւ%q'��������䟎�A�C����vw-�a!� m���-|���4����I� +4^}nJ=��a�QI��{��+��I�*8�`��-��U�dd��F��$$c�,���������uH�L
8�G�o(Z
�z�T���mX���ۙhKҩ)�e�p�K�Y)�f�UZ�BB%�?�jp��sKwȻ��x��h]!T��}���	M3_����(U�3�Ds.)<e-?÷�����P��,��]��k��SO`\f���J�x�:�.�8u���H��!���au}τZ�Tp�Ex�{1͈%5ou�d�y�M޾��x���Q޺��G*�m׽�6h0o��)hN����Q�I��:��;�� J��U�_�i����-U>pl�.Cs�)�~Vu�C�7#��:?f��������5(���1�~54�o
�f{^|#��E@.�y:���b���y��Ɵ!K��2J��L�vط��p�q��֬<�\DK�;��}�N�r�M��P��D���<�Ď�b�;�F�Y)Z{�f�}�y$�ֻ�we��K-7��o*P�7���O(:�*�W������3�-$��ӛ��b�N�A�&V�s.����JC)R�p]6�o���?�Y�Uk|P�����5C-S�(�6��Y�#��&��2�1%yǟRsJm���g#��>�piZ}i|�O��o�S�1
c{s�M�dW��ޖ��	0�7����m(ԫ�E�*�ɮ���vؼހ�kk�ɟ���yfi�mz��5��$���7F ZH�\>���zS��S���[2���B���		�IhX��mCyA�bG��D�;82�<�%8�i��M��5)�z�'`m&��t�ݿ0l�B��p��t���#(�Y�7�e�_��ט
v��VvT��-�N��P^�3��Y�\�jq�a{����[j�>���J��hz�Ɉ�HP)[&1���P�?��⍿-%�l����I4�e���拊5�nc���`rI04M���vPc�r2�L�V��,���[��?e�_���N�k�\�$I�jk*�E�K����i
�0����;t�q�ϔs�q�O�L�����n�8�"�E�GH��˺�W\�̫�6S����C�^��܋���
�����N��a� �OV˺�:�u]�`@��"���G +�/����<��(���CzE%��jk�����2�g�}������H-�P�p7���;dt��]OoE��R�4i8�_87@�Z���̓]�)U߽��Q� �ba24��e��D�D{�?�2m���Ȩ�GK-���£��oނ~y%�LZI��Nq��gۗ$	W_�{=
2�g�}��K���m��*��A�'t���oXv��_F��D�h���-�w���Ĳ������4�R�>K�͞�.c�*q���G�"���q�z�/�W���LB����L�e{D��d���f��,ҡ�9��	��
�h�U��C.�ĺ������[�K�*ۇ��4r3}��RR� Fߛ�##0��/�_Y}�_�;�fV���We9e�^�y�r<6����z�@T1�]D��1�qj[�OI��d���(�1�8[�N�`^X�	�����c]�Y̯��|���ՂQ?*ݯ���͈2�
��d3F7y&걃&l����J@�2T�?4�� q�p4{��TN���l}M��~���[8dW\A�����+e�������!�-)Npxo�c�ὣ��07uc�e�JiOu/	���J���cN�����yXN���P�����X!	���vf�l׍'�I۠�p��6�]���8�֞�B�'g�����2�DeZ^�����-�b�����KFJ�Q$���%�0�xŅ˾�~�"��K�����w�������|�������[-[��a� *c�'i9�=ӯl�\��k�3b'���4WpN6��wP�^�A]�#JӰ�+�׷2�����j�p��v$:Wo�c���_������k>�a�?�#界g�).w�@�Dw����]BI f��2h8hc�1ľ�/�vM���r��"R`a�<�yP
4��$x;�K�G_�n&r
Wڥ���ܰ�}��r��|K��I��c��B�����fX�oc����/\��X�Om䍊Jf�� -�`^��X�Zj�O�=}mF�ϵ�.�q�P]���,��S���:��e���ߒS�ؑ-S�m�wi�,�m,�$�p
|��'L��o�!�!��Z��W�5w�$�.]�v�q[~�����&��kO$��{ �6gu8Vi<N���ۺ�hv�ƥ��v�qwE5LTx���є�ىOrj0L'���'�-�����*�,��w[gҩ�8�l���	�C�Ч*�;nX�R���- FF&o�R���\O���@_WY1��Q������v܃�)q+3q�t�"�ƀ�=����r��P體@��Y������J�FBι"bN2���A��ES-Eu���-�����,oǦ�@5{�V8��+q���N�����G�y[S���FC9�]��UČ��~�5^��z��ݹĤM<�:\�����S8���ƹr���i��P����%��HW����~$�rٰ�>�f����G�A ��@���J�'����5B��AF�j���/�־#HZ���*{�*�nl_	J]�t���̽�ڀ�ǃ�ټ_�b�݅�E��&�»߁��'U ѐ�E�W��o��0X|�\&��h��i1�Yдk�-W5�_+`x�	m0sZ�i��ۖ
�U�1����u!���b�E'�V_�u�b�(�Ԉa�^Kޞ�����@OP���P�lMΝ0A�j���_g�	�eFy,�������_:j�-�4���:�P�+d�;����O�cƎ��(.h�|�ԙ��o�5��:5�)�R~XN.QE=QB~��hxk~�7�b��U\�'��v;��Q���Pח_�d��S6�.g��U�3�P'e�?���Mr%����e*{��
Q���e�#ߣF${<�g��V�g	 �AƆ�����|E�_�'�m�o~�¸E΋���.<[Oڌ���%�C��L��NJ��+��[+��_B�rJwTU��ǣ�����0�x�q��xB,oK����ޚ7ۑ�K�9��5�_9��߲"v�SD����6�W�\`��.�镒���S�� [K�S\��#��[(��`���;����ڏ����YT�F���I��	����m7�I}��9 ��p�i��G���Φ�?�jC8*�K ��8��0��|�t��X�z��d�6�5Tf�$N���9ymL��cht���W��x�M��Gj/��*+{��{wr�����w������S�N�/?��P�>�G&x�ί����:E��ޫ�w�}��s�m�,�3y�a������2ϲEjިh�(SM�ap�h
w� �g��ф[�=����Kc����L�j=	����S��*�`U8�2g�d�C��+��XG�2�~eڡܺ��߻��'�S�(�U��'-�q���4C`��-l,���\ġF�%���kX�b@�@�����綨�P6bY�d��:��F*>�)�1��1����ٙ����"��C�:���x>xB][>�����|e�!|��PG��9V(L ^����i�eU*��B+U�]X2J^I�B�ޛ865R�� �xY4P�my�>�����5�2�YG�o�*�������d���Ο�zR���LE�]"�?��_w��Cg�����^"�<�憺�Υ:]C�cg�����L|���|A�K[��Ɯ���}��+'5�L��]�"�f<��/F��B�T���/m.���w6
�|�*��=���|���v�b�=ia���\
�~���������)j���G����m���b@��M���9�+KJI#���Ul\LzL+oP;��ʆ/�j�Ө����P���8[ 1�O���duf4:�]��c�12hI�F��Q�3�^W���d2� 0CFyC�F(W�Sd&��G�dcuC8U�Q-����i���=�tm	�����I��Q`�B*Q��Vx'y8�	�H�C�Q�p�oir/V��6T��h��#�BA˝�e�x���Z(.a쁲�pI��s�\@����1Ӈ~ <���u����z3+�>$&��z0 A��$����5��D��D�O��Κ_q	�,�̺�F�klB��t%f&(�*��7�lD��X��ᕅ��΂o���~8���'�� e7Q�Z��Sy�A�Sm̺��"K�͚z�|eq�^���% �Ӳ�����p�e�8,V2��gFI[���\��u�i�\`@�s�%K�]=�@�=�Y���,��~�_��l�9�h�u�'2������x(�,�$����
&��!m6�g����6q�K6ɣa&�a��l%�d̛9�<W^�Q��,�mO4�uOĿ�,�jbD�u_��r$cM>�v�?��M?��7��||��˂�$`�JT}z����VFs��\-��^^DW�t-B^߃�՜7�+��itS�`9W���>\�os�]�eS" �qU��01`����q��>�x����VBr��~��.a�+_�\P9Q�U*u��+�1���2�̚ 2L����(3�b�;T]53���?�_\�����a����r7�,ߜ�"����<�Jy�O�O����������6)��R�u�b��i@-�Ԡ�2�=������K=`�[?>�'��[&���H�wjR=Je��^y�U�Ed9ڌ���8�
�����w���nڸ�,��kM^k������I���b�\'�;���"Nybkϳ��j��|Y?���:&�G1�7�f�"�-�a�fW&�'���9�:ćߴ�o��g�P���ҴFמd2J`�J��/���D����J��3�?�fHT��M ��k�����76���!F+���C����HZDwp^tڣ0  ɋ+�ם�J� ��}N]�m}�Fu����u�zK���4��l���<a��;�i����;S�!����K'(�E'�C�%9t�h+���,���I�P������؝�����E�b>Jă�-���9Q�;�s���H� ��N�dMpK]�<U����IJU(�Q_5��H�����\��򏩫�h��f?���YgZr˜��"&�Wx	����k����z�"�jt'X��di��Bq��}��>�z�t��fg<lc���q��+��E.��9p�x���T���m���b%��:���N㻸�e���!:��
��^?�|�l��B�t���j~ ̉��b��M>8��t#���e[�Tituj�]04���#�Y��T@К��9<^����6T���i�siu�u�`��8_tA�Qb"*�m�f/�˒Z����������&�\��I��w��ȩ)���:s�C���;����D��^�M�c��)=�>��t� ��p߶�fx�׏7�vp&��l����Ѧ��SKv[Ga��D�^	�m�1 ��
6K0�:�$�G��P)|���L�HA5P��e,]:���!�R'�c/��X�11*�-Z�������1M7�=*�a��n�lA�

d�C��#`��"^������w->���a���Q�uR�W���w\2�2.�<65��K���40�w��q��ީcӛ���;�#���)Rrf� �Wf9��}���Ӵ`*hf����i��E��M#�k��S\ϰ*�V�.�BGh��zD�e lAe0���1�=��{��2��W�y,;$�bS ŕb��)�2���LQ�l�CB7��vo��^�]�H�QL�qx�J��Cܽq�����}u��)���^2рuQ�P�sp��s��3�m�g�ByɧNQO�r�,���]�]Bm���>� m�#p.~����J׍6U	=%x�9�7
�->j qӕ�����Nf��ɼ�9�\U{z�W�H>�*ZƎh��m��/�tb=ǒʧ�"�p����s�?�gm%�/�>D�
c��h�콬:*�k�o_�J�vIeΨ�J\x��㨖��cCR1�q�h܃�/�&�=��؎�3���,�o�9�^,t��ݗg�E�{��Č	>%4��7�|I���8�������noDdDT��1򩀶��y�� ������8ګ�o�\Ѥ�3T�*�(b�¦P�;������E5J)���"'{��߻���̈�g���Q���=ͻ�Vw���E%MƝ����IUme��ʠ��L���X/�4ehV0]��`�2��~~��e�L�=�L.�&��}��]X$ �z\��~g9��6Ex��y�A�I$���L�����9�mAb��j�/IC�%�ٽ���e� 盃
nc�ռ��ΰnH���F��he��:��M�7Cv/��k�$��(���AN]��ڙ1�c���$����zq�e�[�Bp,;&�ě(���₦�����Ҍ��N���Ɖ�I<0鶍�]~�Ż0II�f���p1�ϥ���&�);��|����?xr�0���PWW���_U�Q��qŉ�1j��0,Z��zA\��9��c��Zwө`�������:#�\��m��$���F����vn����Rȋ8��1b����y;Н@Xq�[RXs�>n� 5�z�%.�!�0@/��3ul���7$��a�m'o&)Q)������f��zt/�����AC�a$KW�O�|U ��:�F�g!$,�>n���kK��FڋL%�P�E<�!��E�L����g<m�ì2q�;d��>�s�5{>)��e�F�Kώ�-m:���em�Ҏ�e��c�p���c�i>g'0��a����u�B��E���/�;�9$00+L�����+��T�X���{g�4>�������/c$n���༱ڬŠ�F��*�@>&x��xKx�~,%km���t�o�������t��h�����}ZO׊�d���7J��U�K�}8�N�hɌ8��Z��j�U�P�*7�:;
�U��sbe*}9�eclf=?Sׅ�*�1�����E(���`�fϠ��l~kI�Ty��̖�S��m]L1���|�K3c8�����M�x�X�e��n�!cs>R�I�]��I,�i�qʅ 6���p@d�!�_�	�6#��ŧ)`8�#+�Mw�Rq��/Jyϧޟ��π$�r�j'�����0=�����c:*{��]_X�|L�"F���h�����,�?ă\�Ѣ�!銥�I�NB������//�~Bﲖ�C�����~��\�1�ƀS�Τ�E}�Z�Ae� �;�����J����p
~�6�,��������H�����]�~{n`��Œ+�R��V��wgaL�Rjn�c- U�73�^��_��^��9�Z�0q�&Z�U���w����Տ4}���z���}hBe8��&�m�X6�bJ*X�5)�|iSdK��bMXT��h@;�֕��	��;BӦy�D̺�Y$M����%�ېԷ�/�+�_Җʀ{SKJ���z��:S?��k�^\���p�� }��@�Ϩ��R�����l]�Fs�p�]H����v��,�/LE�s4�H���7�lĳx����_�˅�
`�_P�B��;n�F���0�
��W����O��8�i�jLY�+?{y�.u$�:R��G'=J�����o�+d�M�~������4;d�=r�b�{���ȫ�Q~�9�6ΙΡF��x��,S��Օ�e5iH��b������f�[����!w/v��,S����K��E)��D��n���a�(T�ߣ���V�=��$޼����K∗�1��U>���ӵ�����#I���q��mBY�(yGZ��/�:0�oL?Y�A$:�ðbJyvW//iY�f#�F���q�P�gs�cc�ɣ�,&�?O���������BJ�k��A�����7�!|��r�	�:��Q���cd�y��)O�I�n����t^|��pg9ܴ6Tq�Yu�N|�E$Hi���,�ፃ��0n (�?3E�"��+//���O ��'1�ȓ��Pzբ�O�5{��a�k��l�_J�X�k���j�#bX3e��V|���<n��mtE�(��	3 0�� 蕠�b�%���7�6��\M2z+��<y�7:s�^ä9�'ݐiV��Lwک�nP
�Yl��L�I1!Y��?��y�Q��+����pg?[�������i�/K��`޽�I�<O�:x��l��rR��)昷�+}�-��#�;ί<֪o�_#�`��
q�D�X`��&�c�O�.̍���擤��򻹠�rk��*�}�W6�RM���M�3�`����v��T�Z�$v�L�H�.�uP׋��"+�a�@��q|�3�tdD&���C�
�j�M�5���	��Tk��s�	va\��`��D���໽0Fd!���3K��� б���PD�ﻀ"�[ENP��|�KͰ&a08������'ٹ���b��2.��g�{��kkJ��u!����>�G�}�X`v_��JY?���nմ�=B(�V5V>�����p�:'�n�9%�Lz/'L��e�x�M#����z
��K*�T���n&�M�ߌ�H�"��%�AM8�+�� ��M�Y�4�����������k~q ������|�9a7I��T���%��P�s&�jP���Q�/,�5Q��P�7��,���M0D*�XKQ+��U&�4Vm�����KaD�۫�q!}�B��Dݳ���U�l��!+����/ĺ�F4�K��>�Z���%������q���U	D��vX
-�=|�q��r�S7�q����cM��_�z ?Q�-Q!�넳�#�:0��q�v,4�v�7��-=��e�g���2�^& V }��k���<�%�Y��}�>�r3��W
�+p��o�
���w�T�(R"�Y��^B����GU��#�r����iZ���nL!��t�/��7|�� {F0����K.:/Wj]R�ʆ������	\����#B��y���b�7���6S�a&�QXI=p�����k<��Mc��*^	n'�p��yCx�@|���?�Q#�`��v�N�W�襙��E����t%�m4�7���D�i�hFv��}}f�ʑ&f���W7&���"��p!�E�vC���V�b������Ғ�3�4o�����Ȍ]c��r�|�uJ�s�>�uK�A��dg�i�$I���W�Pcb �wL����"�ƁB]��=��6J����2ޟ��� ����u�'��K�U���x	�����wۃj�y�c��6f|���e�]MG]�NZ��������"e�K��4H�j6����vO)�V���J�T���$#�r��h���Q�Ģ&���qf|�d!e{�:��q3�`E�i�IB�"���}f�y���AV
rGH}]��_:	i�~�*�ۿzqeB<�e.;�d�����(�����m�������z}Kj�`M�
N���I��npb�C��1;Ț3�I?�Q�����qi��w��'N$�v���f9��B{��qG�,�<%�����]���$����\ж?�
���PE�ceϥ�iH�7`7`���푳{C\KS]Gk�.�$�������j8N岫���)�	�?`+�]��,�̹���Y{�C��!�e�y�\,`�����������ܯ�&�U�j�@����@zk�8�}��6��J�	ȼ�Oj����9	G�'//�u;ȵ�͎��pj���(����ɃAkش4�����N��~�vcxPvm2��Yv����x�+�)��������j����h��O)�1�(�Pǔ�Ьa~b��[����m���g3��J��o��2B1��Brc��у�6���s'�2����+Ӕ�:�?����rd/��'Δ�u����*~8���Ϲ|�5=(k�#����O���	˹oI���m���%�Ƿ]4���[	ӷ�]��D�cjG�1���!Q�tM�B/1jh*&�ms�D�^תIG.$�zM%mjW�oB���B���O��i�,Exhjj��==(���RH�8�r[l�`��2�����o�r���S �����"�0���v}A�I�)��� Y�(�����ώ��v��J]���iI���@i'�
0̅����;�G~k��a.�)=�E�+�sv��-��ο�b�[h�9UD?������D�l�_ُ,a	ڲ�nY��,�W+m�4�7ʕ����$o�5<K�IA""OK	Td$AC������X�ґ���TN̋����"��<�;[1�F��
�Q�P,!48��~�g[�=qB��u�V�`
�g,wW��	�������۔�rn��y��kD8�E�?R>�P��ѻ�U�?4k<l"(3J���w½<�yE"�v��v��"(` �!�噖 =U���6Nz���?�+Σ�1����d��B觲�gV�0-L�%h)e��ɐ�_���x�K�:5,�����2��
���_Fn��0�v����k"�1'�:��^�m����K�!�0\1���jf�jHD|��.�;�����O?u��OE��T�
^���a� ��KV9DVS���	�T��mgo�hߏNJ�߁���"Xg"���y̎�L�=4��+��ի�	Pf�_��:�<�7h@��G$^A�)�(����h�3��	�'��	�s�И�}q�h-�K��}��s���4��8~c�0�?�D&Xȿ�T���C4[�M����A�ө���C�7�i� ���41�`N0Z�h���c��"	�I�y�Ļw���X_����r�j��5�A(F����9��I�9҆^Ģ�eO���8���>��w4_�+[#�޸����$��	�q���FV$�-�
����?������M7��3?�T�0!.ϒ>k]��z�r��g��;��|�3juy��?p�w�fٕkf9FKW3���EG��~l#��O�1}�+e�+�s�]r�J �sc���j����=��и��Ǻ�n��V�&���R?"�2æ�Ql,	��1}'a�ޝ��8q�᝘�=�t���n� x�ms���Us���<�>I�AA].�|��u����ؑ��y��j�(�'�Ϣ�՜�'��.7��ִ�)xW�^����ƺv��)����|6n��s��k��;�P����',3A��U�%�c3E9�1L�+i������dx7�cT4��]���W�us�)�`Cp{L7^%D�PhuH�q�g������Y����k0���x���=�;���_�ȿ8}�HK��!�!�f�`d�=�L#�����D{�(���^���>������qW��O(Hԍ��q�JŞ�Ѿ�!'�X\p�ĳ���u��{4�LQT��;ð�s����R��F��bG�,tO�z%�_T�`�O'k�7�մ�ꗿ���QSu}�;(���ʿV�<��c�X��؈��`���,t�"�*�}�9�;=�фi$#�������@	��GK�ĉW��$ �%��d����-+%0�m��m�RDt�D2ܰ�2�07�FqG��� �
o	7�A~8���ݻ�E�|�a3<�����m���EY��p��*�cܣ6t�j����\0~Hdawt./q�i��e�f��>/d��*�Hp1#0��P�p<���M�>�z [`!!yN��dJ�|@�}���˛O��u�㮇/�
Qy^�F�.�M����|K�A�]�Ez����Va`_��zGxȘm%М�%���-
�`�m�c^��5=�`�6-H�܈�'5�K�H�NM�OsU|%u	u//~���D�|�ql���&o���Z��"��v<�^��$}Rq<O�j_I.����+�WZ� �1�NXKtҲ��4H�'&�����!��ం������0����pɆ�/&����ؒ�Vv2�I�\�D�-sKo��^�Kk���/�@��FP�L���͌b,����4�	h�� �tn��w.uZ]�pl����N�u����ȗƳ����a�)�j����3��(t��$ʙۃ��k��#8�=��K�
~rC�y��U;�]>�����i����%�$;�u�[��4!�'I�����ڋ�#�����˹W�O��?j���X*��M��SC._˃�8)x-<a!�c0��i3i0���c&d����l�ٲY7�e��>���n��k^�5�R��=��r�/e� ����ar�c��n����86v��-��?{�m&,�=vS��ݼ�]���m��0��~��xn f���uA����͞��:��-�Q3��U����Q-��x�d�(�?�j��Q�]�%c�Bc<��ON1X�ê���9�/MS(�C�T�>�skj�_&ϝ-��t���o��"/���"��b$�m@����7��8�	 �42?�\b�@��ɛ�o���ֲ��Ck��^�Z�0b3����?��HJ(&d͎P���h��e%�;]#-�L�i���77����d�F�5��J�߸k��L��G������c�sP�Iͷ(nϐ�Aq$�fH���^�Akz��P�E�YQ*F��3a�'E��;C�� �2�Qv�J�?çx�,O�k�u}�xt��
.�@X�b�ڒߴ���|�����0�]`�k���Ĩ�HVR1ܪ�^�H�{�L��,n���/O�x�Q@b:fu���E��_R�7�~��������
�S�9X Z�>���E)�4y�x5\���?���/��.(� h��_�,�xsam���YF�9(x</���Oǻ�\�
σ�4D��������s�\�5&�䉾���.�Y��܈�ɧp�MA�̸�Y�VY���_e.]���gJl�-xL���u����7�ʂfGv���C�\u:���B;���kXu�W�]��nL6�H#wB_���BA�5]^�h�#�:�,킁�w�B���?b`��H�O���u3�k07���*t���Z�(���F��f��7��=gJȝD���˽�J�A�\lq*��
_��׌(���O%r9���bA�g<�#ʵ�,��֤(��F��x*��j�|��2w�<E���Rܤ.aIeD��>���՜�d��\����Atu������q���i���)���u����R�
� ��z�,7y	��c	+�D'.�%č�!�oWpB��"����֏8�"����"��=�:W"H#����=�\�u0v�_zex��&&(L��Pt��\�>`R�5t���R�C���Ygd�¾���f?d!���3o�Ȁ�(f�ߪ�;1`3`�������/y�4� N�G�[��QV$B
�T����N���h�CI��7��&���kB� �����4��n�d��{k}�G�Q$i?��c�r�w�M��0�(��O�+/�p0u��ꬢ��\����^;�J�U8��>���a�V�����Ś0�u�!��iz�v��۝%H1��G)�J���[9"Sip��.�#?��L���b�骷f*�q��Rcu��7�2��g���PS��T4�����a�b"E��	�H7��eD�dE(�X&�t�Rם��/b@������} Y?���SBNLǠ�x�~Bzh�n���� ,�٫%R7���%/K= j
��Gm�X��M���>��Ǉ��G�s��ܴ٥Ѷ*��/L J�˚����ҒsŖ�F:+��l�h8>
��ޖ�(��[
L�X����^�uRy��˚�S�L8�L��p{�
?�^��e��)�f���.�}<>u
;0��c���n+���oS9cn5��'v[[�Ǎ��w �+�p��\q�2��l�6H�}5������A�.^�ĥ�L� �N�k��CF�l�5x��H���x M�Q��;Ӈ�"]�z�p�w  ϳ�[y��.�u�f���=8�p�i�?]Y�m�򱷸��OK����'4nKa�,��Bo*�C׌͑h��|�<��\��
fՅC	:�_L$Өb��2h�oB���z�7G�h	�Y����4"�\JICo�:���ES�)m;�R<D��� D��	֖:�G�� 7,9��`g̮)�Y�^A�+s��Wa��r�}.�ޅɨ�\\3U��1�j��V����@d��Ŀ����JM/L
�I�v��M��ҙ��k�ikA�J}_3����a7�݅fh����]��c>Y��'Q �����q]�4~�1jε���ne��Ee7'�.eb�P�t�3V��H�Bi�e{lf"��R�k��'��5Na7u�җ��V\���~��]�A&6?��r3�T���@S5���!�0�F}���^U