��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�cޞ���c��v�y�?k	?��m'�67@9%����-RF��g�ϒ���ީ��W��?+ �r��]h/4 �SU����d*�
�����1�d˂�b�V�f�P�(��-{�q��R�8��I�˴E��+RH3�A�`80Vm_�����a�+�oP�$�;�Ț/�7��cg�3�$�)mc�tF��e䬠�՗G}�[���m��D˅K�����3I�w���S���<���#Ya�A�G��|���ǭdF�$��R<W(~-{�l��[8�ʂ�̈́j�m��ԿQ�o�xr#�7*\p�7B�8�K%Z²�FK:�z��5�쁭,��q��@��yH����R6�\�ȸ"߄H�7\�/u��p��Y�J�V8��{ej\��g�
G���|���w����Q�E���(|H�:�]k�h��e<g_$�)�5�KW�/q�|a������� �0��oZ�Qd���=�b/ǆ�C	���l��cq�sʨZ�Np��.�jh��*�X-���'��e�v0�0$Faf�sֵ�y��r2<� [/�m���6�88H�F�y]V�S��Y��Cj`>%f�?�o�BQ����B���F�L�ͬs� �S�3�C#[Or���#;�i7��{����u�^�j�m�Lz�Xt�=�GY7���@au�r��&ö�����F��%���Gx�������Tf$��!��]Y�z^�4�p/J���&����������0;=e^�!�!/(���M����dͶJ�(�<?Q(9ɤ�!�X߇��ؼR��'�p��qp]7�A�����p�dɤ~3�Ĝ��ܘN-%E����\�8ϕo�C'O�����'ϻ��D�^9G ��x�����y�Ԃ�ҾR��J�ڰ"��a�G^4�\/HE���l�Bb$��7$_~BW�ZB_�=�Z;`�Z�fJ�V}܏���+�b�G��V�΍�t*h�=W���������Wݔ	�
9�s9�D��V�-���m�լm0��6}IRbP��kX⊲U6��
{��D�/@ʷ���+�bE��K�~Ww�|�s����#�*?XB��`j�<7����Ӓj)M���q:�v,�4����E��^�!�$&jS*7�l��6g͔I�Na?���eh���ß�v�O4õ8V��6�gg����G\\���ھ&5Vʺz2�����T6�g��$���v�UV�[%Q�+J¯�����x��:��KE��r���>��]���v�?	M�з5��m+�X�6�x��������o~
�=�13l�����4k1A�G�Z�[�g��_:�k�#<�\�0�v4_����Y^��=��:�[w@�k��xH��jJ�h
3�޼��js4�qWȚ^W�J�1[���Y7��Tc�4 ������������{�]���ٖ�i�^&�j��	��{�QX��Ѥ�j/��/��D�p��S6�2�q�1�j����6� ��0>����QR]rGb���~�҃
Яq�e������!����K5�!˦�P�\�"s���N��[�oN@��;�� 何/f &����G�@�4V��C�-N���~L����M�IE#�S_�iu��D��]�a�J=�����:m����2�@��'�;%͆��kp؉y�$���;W�a Xhl��J{`5`���3S��_K��O�ΪX�\��&,��c&X�Ū���y��o��B��H��S���r�ᚷ�|1{P>�`�P�������v�e	}T���d���+��6}�m:f�&Ռ!�8�[E�\렠�(X!�9k��%�W��]]#�S��UR�#/�}�i\ɺ��{��Xܺ�2�i}��7K<|����K�2����#K��R�����f0(�����>��RuC�~��]��${֥��|��;��kjm��m��<��s�Sm�+ӑ�JSNH�+)\�wW��}��Y���-d0F��z�s��P����㤵)!���Iyz�[�������r��;��\a�`Dfw���E��di�d˛���H��ѳƯ&����J�'�q��3�R�u�4��#1ؗ�X3-zbŕ��>^��`�P�U�OAk�P)��7P9y��_����8F�8el�7�b�{�t��
r��|����pK��]\",/�Hԁ�����
ѡ�B̙Z�L���4�c:
�0g�.E��_N�>ܹ�!a�Q}L��4?#{Q�	��'ݱvM�P��TE�n��l뮋�^=�G�t�ku��~Y�9|����)_~ӧ��������o�a�`r��Ɛ5���'u�x}��~?5$9�"/R-�n����ub
�U������ε6D��09�ʂ����B�/���0f��
�kQj�Q�j�-q����<N�6{��/f
`�P��g)����r�腤ڰ�	+<��MsbM�̈́��b��.CF�/LBkI��K1:�^�/���"����f�)bF��ujtzLd36�?�3�?�\����:�G�����rˠ �}%�'*?�2�r
yWP2�Dܗ�ۛ0uRE/ն�=V0a�0U}h�	G�$��
gH�<�%XUL�0� ��݄`cR8?�,�['F�~:���� B����Ӹ��:������E�h��'C�f$2�k��h�cH\��|�$���t���(�>8$�#�1����Ǻ�fk�¤��Ü4�/EA9���\�3�6�8Y낵�ܛ�VS�~Y��  ؿ��(����M��u1�]�=�D��Db)�{���wy�簼v���&��� �a�K$yYΥ���D��,�?@����eU2���o�Q�q�m<4�X�ԍ
�����n��L嚯ֱ��^
��v�vE�o�F�L�+�ꑭ�:�cY�HN����w.�}����}7��4ap�m��_Z^w��怰�"(١�l���g�� ���U%��6(�>'� Жl]�{���X ���w�8�J�3fQK�Ή������]�3��/�K�o#9���$��9^�n�̱�@iϼPd�����3�U�H:Nۈ��E/� �/t��k�j�7߳3�����2ĩ�8�g��dɓ����C!�z��:��΢-"����(c�� �D6���d�q�b׼|MN5$���;l�	�w9���ސJ��.�/�q��������J��j��B�~�|���+%?N�,�wQ&�D̅�U�?啫�)�VN�\!�q�?�3��*-�͑b�u�~4����?�	d7�X������;�����k0���67��o�߿*�Ɗ�%3��W�T�k��ƛ������Ƞ(��!�`�ÊZ��Rt�����H��|9x5w� v�sj�;��TuBs�~G�z��<2K����������%���&݉Z�h[��V��S��.�Ǉ��g�~��=6�/ ?4��|��{Ң���	0BZ���|miI�I� ���-yК�\b�?�;��4���C8�ti�zh���G)Y��?}�HD^2��G��o�[��y�<�.tu�T��_	�Fa|��?T1/�rt.`�^�J���c�)}XN��}l�ŝ����t+_��x���bG���9���9|Ր��?�3o�J�#��TbS��)���3Q�V�1�
!�:q41��ʊ��g��C�U��i=.j��s;֍$=�Sp_M@��_(�!̅�ۙ��EߚS)�}�0�7k�ڈP�,���wI~�| Mq}�RD�8"���,�&y4�G�TAK��J�����_&!���\�^&*��B�lVڝ�\J4	�e#��A�� ��t��`/⏕`h(C���ED��m\�?����P;�|��HM\���ܵ�F`F��%�4�x[��kczC�	1�GνN�H �O5���|Z�
D�i�4Px��|����?c8���:�m�^�ԅ�j��D��cz���qI��5�����(<	F-~����7��f�(���r�݂��:�a'�-�$`jO�M� �:O(��-�\���o�,m�m�vj�M�3�/�槇��4���?�������Epg,�ٽ������d���esl�����h����������b�f�����9l��4��Zz����X
����2��CDy���X��xOY�a�����UZ�E'�u��fy6��'��BOď��C�6Z��Ѫ�xf94$I+����_��+��о��"Op��t�d���@a�ky�A��x��ܨ�}�Ώ
6M.�O����!�G|���h�i������e�F�=)^��zIW��c�����m��hF�JK��S�P�;؞��x��G�wb�?/
����F��g��2/ΧђO�Γ>���\�HV�I�/]�ȶ\o�F�r�S��x =�k�h,B��.�B��|�.(��ŷ� X�X�Ĭ��s<��PI2���D�;����K�w�2q����XW�wIm,n��q�7���E���m˒��i����79¨8wuM$�����8�YR��R�1��_1OF�B� ���=�W��b�seJ��.�T�#P��3$l]����W�b�2���gn�!�mD��HL���|��T�̶aO{9�q��<�p�ۊ}9�QQ���3���eP���#vz~l�O��H�.��.��xւ�8�;A���X�'m�SI�K�y�Ӷ�_�}ڈi�QX[�(�J���7C�!ΠC�k��ޅ|\���Asht�e!�zxJ\�|>��h5)8w1�k��D�ҟ?t�:RtM�����F�tYՖ��Phm���:h�(6ͤK�۞m��,i�
x�Fv` jP�;�C/���d�r�䬪E���JX>��`~1��Ya`��@���<Q�=�г�y�A����P�?Ξ���E�Z-!��e��kIy��P���'���x28�p"�u�$��ٲϮغ��*;�>��
$<K������0Щ�B���"�@ o>y��Y���Y���뱐�LJ�jKǛ����fu�5c$�e�������?8���do�}�Z`'x>%�C=��
�bEy�t��g D�F�8OL�O�׌{�-�������Z���
�5�E��.���q�(��tN�|c�X|x	���s�5�Ԥl�U8"3s���e�� �g	�ҁ�N�~�X�W��:ٲsY(������5l2�ġ��;ԑ*�V˜�IY�&��cEpN��7<a�s-�Z$P-�ϧ��<V˧|U�xIz��5☩R)9ad~�Pv��=U�"��7E��OyÊ%�}�U��	����ǖ��;X®��@�0&�����}�_v�K����Y�M�a��?=���V#_�_�[�����iiQ�~@J�^����l좙K�CSDҙi��������o�ߊ�hB�UX5��*���m���Y����Ôn�Aֵ�� {�܂��4�	���Z�r�[s��s[[%G�9�p�����V[���s���Z��n�x��qb�o�x[����[�+�B�),�g#��u�S�.�P��Ǒ���]'��E��pc��؉&cy{�����e�4���5���� ���4����/3�~j�  %�<��������B���񰲆��y�C!�~���1ȕ�,�0n?��-5�!P:���KL�{�k~���t������i���~�����1 rpa���#�W$K	mm�x�;V%�p|%w��?o�eq�e�����)ɢ[����j_����9�BU��ׯ��9D�͏�3�ws�طe�iԹ]c���,x��܂����U)�����9֊��w�s��	`�[���	�B���8+��J��|�Aь�ѧ�ƺ3�A��&H�Kq�b�{��:#�Z�7�BR>PaLr�n�f��D��]�ՙ?�������ؗ��x�gmT�/�,�v�m�.L.Ka�����6�zo���@��?E���LO�)���^�z4��F�r������E�o�'w�F��ZEF�9�/K*7�^�.�C���m�${[����8��>+h˅;!pf�sj����] �Y�����e��5��+Mt�/G���9s��n�""�(�V�L�^�{\d`U�A%��E>@����w���6�Y�"����!���7<���S�t�{bc��}�~+z��`�&��O�C�dxdD�QT5��7�iܲݍ34��h��ƉQ=%�����(c�(� Bl:s������Z>΢��bI�9ԇ���$	�����Q�9 f���zLsA���q����A-f�fBI"� ȍ!�m�r9.�z��͂�F����y�&����7�LH��*=��d!o�4�2<���~>^7+ښ��G�@e����B?�Yb05��Y�(B,�UEz�J+�������@K��1�~��I������^���/FST!����`�__~()�=nL���e�(Nۯ��6�[/��mKS�é���B�� ���_5��N�v,�j�������U=5��O�"~��S=�B;����f��j���{���e�G,N�Yސ~gv���Wc�xP��:�������&��ud������x�ER��PG��ݲi�f���y:�c����������0j?��A�7\���Jbp%5Tlj�
[�0�]`�R?��4�g��JE��<%����f�� ���)N�H�@������L@���{/��أ�O�ۡN[��oHE)O�a�����}��k6u��Q !��CL:�cb����J�4� ����.��c�'kf��s�YśXf�S75��]4$�F^i���k�,a�����O�s/w��+�NS
*��c賤�<N�ֽ]�Q��eCw�=�m,��[�؂�U+L�y�غu��s_���i�HI����z���mZ�U�1q��P���{5�*p�i�	�j/!SJ�� >G���}&~�f�,�C�s���s���)cMϺ
�guz�i�r��Ӭ����2�J)�P?*z��A�-m>�������L�����upy�`�X��
}ӿ�[>�rm���V��`�|�Cp#�f��bvB=_�;�.븇��J�q��e�k\G��k�t$:|�af����5��5=�����U"Ϟ`	�������ύ�, j~�7iGlQ�� ��p^�r�3W�:W=[FܒXF����"Кdk��?B\p���g���4�ߜ�@#��χr��|nSd�\�\E��.����2}��P�v_�|4�.�5ڈ%^�������5�9��л��E������*Be��[�.̞��/�,�3BsO��/w��<b�lK  p�P�x깕�	#��%i�h��T7����T�����q$ѭ{��_v���
���ke NÓ�?�!S�v��s'Xz�
�6ܟ�L�E�)���N�H_�%;1�A��&2�w#O)�%�ߓ�>珃�Ҙ��H[�w��w�ċq������{�!��Gd���N�j����(��?�&m$Z'�T贝�SQs�_�=!��d�9�.n	���=9Ҫ����Z&|���fG �Y��)���Li��V�1�P��(�%5�`җ�my���b��7�k�\���o�U�k�7n�y���8����f�Ē$`̦��ˢ �3�"�dN�C5���+��C�J=�i�I��vX �whW�൏�H�Rһ�0{�Șe9ڏ�O�6�д�B!��ԇ��#��S&-��o�X��
>0�_k`w���s��NC] �����5���Ƞ��j�k)�7��-p�p���J�����<���+#�\O죝3{}('������8�E��4�ĉ.l��X��I;~�
�\�Q�f
�謃;�K��0�n@y%R��,6cf�h�����z^A���`��0��룱Q�ћoQ9�?�Y'7xi�� ���EǝSP��?���s��G�Qݷ���l#���WQ�
��+>�K�ž�X���=b�m����$��7�� ��p�T9@(�n� �!&N��
.I�ٱ�����U|A{m�ѥ�V�wU%+�[�.�μ~Aq������>E[g�}��T��s�[���ŭN+�I����V�m�
��mM�V1 ����WS)]_���2��b�$�$s��(�SA4��s�D�c��3��� ��B=j*�I#f��c���-���;�I���*�#��)� ��,���EF68T��=Na�S@a5� 50&kCm���3}mߙN���)���ܶ9���j��e��h���������>��T��l�2Yќ_i�)��[���I���Ŭ�ّb��iTspc��)~�D�z�$�UĽh�S�������ے8MV�V�~��d!uN2�-�f�^��-��*��� ���(>0|��+�O*�2����N�I�!�/&�ʫ����~����A�7^A�ܖCUsPWR��\v�΋j�]/����`%��S�x���m�9�_�2�D��ث`U�^�ꩃ�c�a���J��#]����'���蓮��~x��%�)=
�Q��������>�a
ٗ7�dr��ƌ)�8s��Ė|Q��Îd��>��@d8�������7⻒Ia��=��f}�Q=��]���+tL�,��'��)Ci!�~���r^���Δ��2��X� �QfiQ����d�G�n�s��p�;��2�+���}��W"��d���aC��2��V�H5�;!�K�lz���-J-������	W��Ès5�{��<�_�"�2��o���F�i�w��|�!b��Zs�`���~��E��d�Pp��s��Yη�#��f�Q`[JK7ќR�ݏ�Qy�ac�(�)��%F˿\��t7���7��6��B\g��`�r��cY���
��#_)�b\D޷ V�熅)<�E�裙ቜ�3w6�y\����N������y4�]��Qi�U.�/�^���v��^4�W%z�L�1)ğ��'�唥;���x��b!ju{�~�ah���5w�$�qnݞ��s�x�y";|�T��8�b�EҲq��h�ng����a.h��/����)��W'��q����=�����P��+�MӶ
^�#�G)`G����b��D���M�x;)�������$�X�DiW�n���C���\���}�v��r���[۬8+i�9䠻l�n�2I�\N.�)|�I�l-X���:���	?}���8�]z���UC_��}V�L��o��a�Lp����8��5����w
�f�ϪI"��U�|f9���[۝�g��v������kvk��ζ�sbq�U�F܇RjSI��T����vv}c�GwP��*#�)���pg��65��&��[�ܬ>+��`����$�d�����N&�I�Ԥ H,�6�s��	ϻ�7�w;�q�'�����dX@*t;q/z�.�sz��N�����e�NX)��Is�~uKؙ\��������l�yW<���;gL�)e1��q�\�c�xY#����<t�{��j�H�����͇?�W��Z��R�]�������'���X���π������1��e ��+�÷�Q!Hぐ��z��5�&g��#Z�����U�&#f������jg�B�]���B�(O������D��eo�Ҟi˸��49�n�9j�6�i���Ł
бXyϯe�ȷ��p�+m��Gz���������+���=�@�i8� 1G[��_�"�QC8� I���;rUݔ�D�	���M∄�@J@!3�e���6)���"�����t�kH��Je'���KF�����9鍯߷�R�l#҄��Ŭ�{�wg0l��K��$(������g�O�=�� ]=-W�r}t�k�G �	N�i('g��7U���
���s]��ND��QεI0��\gUJq!nHs]T�$Aj��_�� 纣 =<��q͞�"��~����I+��'��f�O��a$�"�#�7���|Y��=j8b��5�z�<�3�J����-N;�����vJO���+�R������Hs��"t��7Bc�B��7<ƶ4��Ǿ-�Sgא��3���ڒ�<��\;(�z�vt��I���^��2��Lb8!p2y���y<uƩ��wx-y�1��0�$������\�}�.���`z�}c]4������]�ГAP/!B_*�N�T��0��L�����6~���X	�	'0���?N�u���0����K� �e�v�䱪ˉ��*�>�\��-+$^����f[X��o�#w`�@��� B�F��+9���6�{�!�������˕���K�<=�)�5PeJ�����Jɍek�[}U�m��{?@�K�YGUXn����)9&�|�h��~<��cw��j�vM���c���H��m�_0��Q�����Ƣ�c�W���;F]{^�M_�O���A6�������(���n�]�<��2`"��_�od�]��jI�B�R5y����mbv�k���УU�ͩH�eZWg���` ���׮q����4���	 ��_��O2��䴫mD=��kk&�����mk���tu����O���!���m!P�Q��'��	%���Lb��Jbc�[F�Ho�e`��W�,�e>W_����hЊ��PfV`�Z�TF̰a`��ȣ�)�P4!l���O)�
D���cf���q3h����3v��PQ��Q��2u�e��#�����ѷ[�����yr�����PQ��w�w�R=ӿa�>�u����{$5��W��|zǸ�Hs�#�E�qo.��x�E6��Z��+pL���
0�1I�F��2N#�����vFT	�T�ᗽ��;�?��a�Ȅ~�^�HHo��d}�tƐ1�`��&i�IQsiI[|��j*՜Ļ����(y�vxdp�آ�G hw_�|�����'%�v�������pv�(�{9�z��_��m��-S�Zú��`�Zj�#S��WMv��S���Ü��T���K���.p3C��e|�ר�C[)|ŏ�	�sy�ܣ�)�Z��
�A;rp��r}eNk**T�~��Zl�Xvl	žj�+cѨ��K'Tm�:ƹ���yj�]�����A�P5c4)�F����Ѓ{�H��L'��l��3���������vV�\) �pȇ`J�
�R'�9/6Ԥ-V���Aʥ�Я�	�pON�Ɠ���'�2&��~|��#!�<��Հ)�!��䚲{\ӠS5�Xky��0��*������ybq�&,��b�%^��b0�N���l�@5����m�Rǋ�f�+=�`�ٿ�p�&���f�˼��s����Xb�O��B��M�l�)�庩
�`
=�����b��I7���jbR�z=(��C¾B.	j��W��]�$ɦ=%�>�g��^w[/�H,y#c�ߜ����̡�z�&��/0|�M�(��)v
\w��Ԁ����,�<Tf@ޘ��1��h�M�
�!.���Þ�����n��'�9��V�S���ۡ��kU���&_��y,ml�l��Y��%>�^9�?F^��/�5�"
U�о7=lR_/ �r��N&���d����u;�Aޘ��^�W��F����+�����o�Z60��4ڼ��J�%2����L#!DH��3_��@��&�#�h�����D2�0�p�,	2:�@ �El����K�9i7�Ɗ��ڰ�a�ꍚ�B�3w`���!`~�B��!���A��2-���T�A���V�~�)�V�R`��|nSz�-ϟ��lYI��-X�$��j��A �)9K�=��,���C/�t=���Qq�G}#s나�c�=x6���Bk1�r]d��4�Ɖ�3*؄)4�~pMM:_Q�������,-��eI�x��[j�e<�)��?t�ӟV�Ʈ��� ��q8l��䔅g��u�����P���r��ޟzwut��.�Q�s���,�zC�VP�t�sR�sERo�_���j��f`��ĝ�?�|�J��e�eZ�Ί�~��7�a�e��<ܱ�p�P$��\EK¤-��,F��H`# ��]�п��7�m�� ֹ�����`��֛L�m뿬�)Ns�Q`�E�l���H����'�+�e_v$�C��z���G/���v$l9��nL�Z��Sqlo��~�R�$���{�c�ƶOkx�gyOďji��ēC�_*��"���d*g�D�!v�E��za��m��_(y��;Z�����3�b�~�M�۞"�wْ� ��.!yF����9�mV_7��z��_'f�9�������ǽJH�ˊlX'��o��d#1|�)��!H�ʽ�x1�Q�/�$؏��6��qhl\]/��&K��Q�ֳ%���ݚ/��i���(Zx�t`�C^3��Z�I�Tl��U^��;/��v3�����1��o�1>F���./j�
 �^2R��~L��y��R'��?AD˻��ߏ��s���@�Vf���`7�,]�Ii2���tD�"�1��~�0�z@h�0���]2���JЕ@:oU�욮_W�U��S���Z�[?$(ѵ;۶���SuZ,�#B�<�cA�| �1�Ud�	�|��q`���Z���7� エ��E�5V����J s
��w[w��#e��qd��f���p���e�A����{����R���^��4L��naMN�[]/��+�4�n�}�Y*4���r�̞h�����Hk-�To��G����LQ3�;�)H��S�+�x��;�2��\�-�-�"�2d�U�e�~Q ��n�fkz��Hz�N�x;�Ӿ)O�D��a��B��}�d�O;R��������p�,TO�����RO3�4C��	3]d3gE&���P��#cHp����׊$SF�>���wWUܯX��ץ��Y.�8��[����������u�T%���$?I�y�?�`��B���#��yP�S����Q��ɕ\�;��0y�+�u<�GP��,� r\jC".Y�e�4������@72|���[��qQCYɄvaQ�u������\1���>q������.�YY����KS.3^�=����!�� ��`����sE�u��ܵa�i����7���ǖi۪UD��:���I"�+k�ւ�~�G� nޭp&���q��$����X�PY����X��H��4?1SP(�UY_��F_Lq�?!�Ԉ�������}�WK#�����ql,`.N ��r���+�;��;��vW�m����������&j\X����{
�	��gk����!��h�s\��츨�l�x1��b ��[Bpz���@s��һC�9?T䳙�ҝ�o+#q��$#[� =�z`��V]���	{��@�X�]>�R6Z�t~�;��/��v���{�R��75���H!�@�5�������!O�(2I�"^��z���E�ز��W�[�Е���!�<�� �e�E�gǿ���P��4�Kh�6T;H��"Eu"T��
H�~(Q*�aLB�eacs�6�0}&��C�o�
���s~n( ��B�+Mg��k���{��kOu;2�9��	��*O]x.�'�צ�K	��� 5�I�+��}�f���������2p�M�E&A�|X��] �C���Z����W�⦳f����yζ���b�6�0vп�F��$�`ӕ#rNG�2����WF�O+��/�(n,�.�$S�8�q���˦&���7|E�Z�?-M�G���H�v��>Ty
X\(��[<�kH�生��ם7BH�+�P>�1?��$��*s�YلZ��Y�Ɗ^��v�ky��G�_=�����1�{W%VG������`8�J�H�<U(`	+?���L6��7���|vD:;u���P\/l�l�C��U"I�^bk��uJ%�z
~��v�ؘ�ݱAA�'��P��h�-��O/S�+|�� ��Mi��$��B�������9/���ͼ� e_p��CSe8�w���X����%�r�m�2�>��˚���PrW<�W��-����`O�}�<�C2��ți>��:�q�Q������N�؄g����S���\��+!���<��j��R
+��$ �V��0�0j�*	�W�h�).��0qc�V� �tR �rם�p���C�] �^7$Y,��z�y�
�m �U�����G�((f>H�x�N��#�Z}���:o�.o�t?x��kf�_N߹��5P�� }��uw�&~7I/d��|�z%&!����:<����������k�����\�qX�!�|e�F�un��{���U�$�����r/2�J�U-��f�	}Ԭ	���큧�y�yㄸ����-�K�\&'`���n�����Xg-��&�-ߕ������"�f�*�s=Bb[;�N/��w�)�C(��+^k/�yر`/F���M�ֲ�%���I�F�:F�����A�+O���T�m�?��у����p�������Qj���ʹ�q��)y�z�}�rm(�dЖ3�T��|�b'�-F�XmCy����TY��3�~�z��H�Tg�6I:1���]C�R>v���<���e(�����0��ċϴ��C�qZ�m�H�{��k�mSBY�O���vn�y:��� aF�T��ZŰc�t��H�����&8{K��d}���*�sAХ���(�g��1*�v4~��t���1C�"���=�����Ѵ�v?�*��SK��l9�l�r��ouv٦/M���&�[�W)��5߼�1l����҉sY=<�;v8P��<���8�����
��̃-������ݷ<7rKc��	�I�F�h/���f�N��o�.��PWD�ʖ$ؿij,��F�n�������������K�yL�(���e�����ݚU${ʲ�"i&�!ibu���p�A%3c�"k��0q¯� �r_�x����$�=�  m�L����fܒ�CoDJ�@��X2�O��N�RVՔ�*���jZ��@��v����7�� t�3�����?T�#�z���ĥH<̕s������Q�����Sz�#l\ÎB�P�F�x��%l���F���jv�?�uH1�Wl�'e��sX��
�d�}8@$1����t�N���7W��k��#�������0�S�v��%B��q������l�ҠH(�#h���P�Rtn��m,�6l��XP�_)jv+��Ui|��-�z@�B��~���6]C1�����<�|)��w�<$�¥��ӌ<����R9��]B��%��/��js-n�� {�Δ�4���a�f$������j�n��}��<Q
o��d�\[��K.�J�F�X2uD��������u0̸�b�K�%>�4�?�������Np�Yۅ����ȇuc�wc�hΏ���,�12(c?�OMyUw��ԧ��H�p0��3a\RA�^�-���	�uenO�[��q2�$�cm�9���\)\r��z��ƴԔT�9�:�U	��06,�:�Ӝ^J��w¯�Kg��eз�_���8Јڮ�u�j�༌������gZ>6��������4�N�4��l��3s�t���8��i)Y�]����Q<���K@��Z�8lsX;�uT� ���c���k�>=5�P�T]i�<zH���
�]�1����3�D������L�s���|�B}����噎`��4	��C9
�@[: �D�ړ�`�<@ɘ�qʮ�IXFؑ��F��Je[�Ji�F�`�z\�{Y���_�·�h�m��rp��QQ���[����tqbD��I6Z2�����x�ߺ����}<}TI�$Y��*b:�m0��h/E��>����:0DFf��!ߋӡ�n%�7�� e��|ǘ �SA� ��}�l�`D&= T%Д.��]���P����b��p�:]�aS^*���M��37�����2>�x�b��)s�PD+�Nm�_��A�*�IH�3��ڮQ�p'�K�QL��Y���25O�[� %��`&�N�_�'���rߠ�����5.��눀��^��
��:#������=4LKg�Mup�� ��<<m+0�����gE	P*b����#:Y��|��o��;��#��2�@K�.�6Y���#zȺ�6���3����?����t�5����|����uXDlU�/�oX�-���{H��^d�X>!!-pL�w��onk�}w���[i�x<	���I�t�j��z�O�*܁=ēd4H�@�_�"���T^'��fm�Wb�#���\T�%�t(����P�k]!:|��|J4���"�>f=��"����i#+��)@~��.�{{�l�F!a��e������{��̖����O���0�M,H�')�ޖx�Y������*з��x�)�nE\5Εv�h#��a
��}3����Қ.��W���Y�;�i:nա�`y�-v�8���F���\3�Ɖ���%/M��%�dF[�3���=H�wb�1M,mU4d��G�i�/m%��?1���7QM�e
��`;8�ţDO���@)���;��R�t��n�Iƥ5z���6yZ������_=�f����u�̞b�i=�O�eH�� �<X	�h-�$�y�9e�Y�
��K�M�n�mZγ1+�P��
`6�0�s\�_����,p�T1��:��\ިw�R�cA�Ax�\����˰l�	��X��H�g�������߱b�<$���VZ>G���V$|~���V��r�,@��{)[A|u�Y��#;9~�&��Ս�d����L�#3�iF� �gcv_i�%e��+7	ff�w���Yձ�����z�D��F���$���P��#ϥPHyo�18:
��
Ϊ�l�dU�7PR�i"U��7�Ԙ�X7n?X������U�>)�C"����M�9.4���7��m�������q7����X(t��A5"�������r뙾�=Ҿc�i�.d�ҷMs�I����D��-^��%�ͮ�[�x�c��lZ�c�ES D�$0ޣ�����R��&*���y\��T��j���"p-��O��}ҟG	~��p���Os_���S���l�*+�hVrS�����׹r  ���R��T��ã[c)D5-�D�]2��i?[�>��qLS�M>r��2���0� ��@�=�ˤ�j�� ���ZZ\D���T����R���oxd�r6��c��3��0�&�#��@��mJ]f�w�[�k�
��b�!���r�D����b��$��p���ڌ��@@ )9;����ۓe�nmjP��L����/�p�<��%�P$��{���1�����h�xyq� ��)�,u"�"�;�3b��?א]�����I��%>�4a��Ęf��!��<� �?C��b�+D�h�īW�\`̰��v?�y�-�k�����Rr����(Z���FC��������5^匕^.K2b:�o2�z�ִ�_�͔��9��X���!�5�`�Ւ�u��؜Ă���O#���� m-٨����1p�p��t���/G�c�E�	���y�Pn0�^�+��	p����D�NZ�����ߓ�Zͫ��ɻ��H�"�g*bK�+8��b8�r�"!��|�P��I?����A�{	L��lf�傕%ޏ�8OZї�>K>lƫ�[;N��1���M�m�c(�`�o<�������u|1��� d.�X���0r�s>���O��!ǣ�V��b��u��9�%v�?;}����Ӟ�n�j��xͼr�U�H��1��gsE��߿䌩 E4��8�8,��@.���2�׍6p��o	�rNZ��4�7�^4f��
�!�.��|E*E�-�XHG�q	q�@D1����	�]��r��{�bЊT��̐~�T�>-7�� �6����[]<��q��K�㢩+�����Nx��#�-k�%��~Q�8l�FWޙ*����9����|��E*���t���J4�}�n���1�8�_�)\R=,6]������>��d�J#t"����X��Fb�On�]�!�^�*����o]�$�x��L֪i��j��0R=��]Ы}o�\?�z٠va_���C7�T��̰�����܌��&�*7%L���i�Q[���/����𖯙hZ�������w��f�R�aV��\|6�+�>�Lc�˯l��=���Ckb�AA�!��b�7��w3�7��P�>n��xF�cy��Ʃ��K�e����կ�- ��!qu���8�x!C�Yӟ�%�WX�b��e��'q��p���jU;[�u�fl>GuD�J~	i����\�l]-�:�(f~�&��1ٙpǹ�Z}NqO\O!(S�V���L�����F0��`!k�9Wv��@:1�C�;_<cot�TOHh��~}%�M�ߤ�w��ƫ�.�pY.��%3�̼L������"����ޚ��1 �t��� �組M$:aZxH�P�ݎMᦨ�����0@u�-��I�r�mm���I�����@��RZi�(�! ��+d:�����?��]�7�3�B!=�9'Kj���nTy�����?���~;j�����3��)�1����a��y{C@��[�g�2;�<�{0%��qs/ e�<7����J¿!��D������c��Fi= �G�=��t��Q��*]z�a%-�����?���2U{���O���	m���	�K
{z�ťJ=^�'�g�w
�u�xw��Y�U��@F(HA݋`��s<����mщ�,��j��R�n��(\F�6��Vl�����{�� ��(R�'%��_!��9���~t��5�?0�l���GTk�NJ��N�x#Z�3lђ��mq���a�1j��"p֫dqC��W�T��F��ա�mqv� l�lՇ���"�Ӭs��+����%v�6���n޵O�[��;�-��5��γv�F�>��rcan�Uǁw�_?bJ�!FH���v�:$٦څtۖ�J����cpM�����-�lsj��n6��CQ�NujÝ��wqZ&7�;)bw�{�+��^#���B�� ����nE��zW���Rz�fJ@���U2���`Qk�+}�Y��D����R�l>�O!����m�Iܢ�Ղ�)���}�O&M�u@9<D�l�\�1Z��q�#̈́�t��e�t�k�xn��Ԅ��8�|�u__\!lfj��8V+H���C����,�D������}q�$�=�[�ò��#�̂�|�C��$��� ��D��ôК�#6�+KΈ�7��k)uh�'��2U9���Q7Ŕ�4��gv������5W�o2+Y�p�`W�n�W2���,�ʎ��_6X�y�g�=h�7����غ���xOd��i�+�\����V�fK����AR;a��J�o�v�)ܺ�'�X�W^Ͱ7������\ϿݱS񳿉aVK�������s�1Y�X��l�����=�����P�&���aBh��I���A����Ԝwډ��� ��@�E�\q�-��TN)�뫧��◈�����؋L�%��"�TaF�P"2Vfo�x=��1{���$g����<x`��7�.��Z�Ⱦ����J�$��{G��f���T6`�Â|\��m�BnodnW�	=Gj�ă�o�F��N�H�$�Z,��C3���:g?hJ�@3�s/����z��*�6����X��j�[o$ϳk�4�։ư+^6t�i���r~Mkkp��@�&�0��*|�]�(ׯ�ƦᅪL�p>�4
F��3���ԑ�45����o����/�<��P"[���!0��|bES���UAH/�/�㨫z5m�/��W�!�����cr,
���n�!�z���aqUB���5����N��,��)���&�([�kڬe�{�S�g2ZP��s!��2"ֽ��C�l=Z�Y�T|��8���i������w���A�`��P�9�������eo�rQ���}�hW�|���Ӏv��Q]A=�
5�UHBC`/HP˦��7�����k�a�Vu�p����������C���`_�U�í����m��]|+�?<�_��̍���A��g
����U�F���"޺x�$�W�~�#����W�z����>E�.���J��]P�Ѝ�%�L7�/$�\�'��s����-(RU|���9�ă�l���':0�4b�%�⯫��#��,e�0��J�בd'狙�?gy�7]}�!A�=n�{Cψ�����E����`%"=�~���5C���
b��>˙u
��M<�t/lX��D7O�yY&��"Y6턓�ڇd���X{�TU���U�����N�q�1|h����_�G*�d�j�L
�X���Ȁ?D�`����`����P��Ӌ�����2����n���L���u��[v�i*�'C��`d��8-/g�ϰx�ڔg�����s��%�D��P_J)02&մ�����|eB��ڙ�1�6��v�$�n�#ߐ=��DlÀ��?A�*��u��epnJ���)���4�I�Vܘ�˝~��bA�<��_Q�Ae����lP�S��Zk��ϋ�n	�O���O��Ũn@�g���F�l��w섉ۑ#t;1e��v��0}3�*������*C5$#0D����0]��W+�7�F=��m�ķj�:\�!Ei@�鞳��j��Ȉ���``�V�G"�ѱFuGvSo��$svyP�M���$owhK������VH�������J�� 9ޏ�����-`�.9�
+t8����c8����GmR���zQ�C����	�u�u���UDI��{'��_��=��]�y��;E�%CX��j8��`��S��jٲ��>�ɯuTN���v��4��q&s{u^T<$zH6��I5^<��*R���TKB�7h���tx
�2�*��y��W$�wj�E��M�T@��N�B=zW�Z�������9�`���	qO�L�3u����?���S����pR�=f����!�i܅�er+긙�߰4�m��id�?I;@On�S���Ⱦ��ŗ��e�+�+�0�o�b�pPvpЀ6��0gb=� iM�	s�&q�t�ԟ�&V`��;����}W�hZ�4L�������ԏ�+蠂�`[�M1	�����M�B����=�Ǉl��Q����=%e��χ�L<�e~��U㭪�������-z��j��"L�N��|0�� [����O�'�A��p���7��ܟ`���B8x���"�X�^5r� ���4͎��b�) r�X�F(��*�g�~��Fj
�_�0�����$�@p���؍S�� �#��}D�Mԫ�g#{�񂂪���ɉ��F��$c����L�:�Foם�S�CcE:�#9!h�Tp��墸y/��μ�����#����c�I|3��]�o`������q�J����q,�̚%�T�if{��H#�B��4`���A�6)��J�T�Y����9�hyġI$޿�ҵp|n��δ�z�2�����=���<?�����p j���|�|��3���NՎ�q�_����w�UV��<K4�q=��XgVjh*��d� ��)F�@���>)I��<y_Ā����,��0�(ç�8)��_�.O�"%���)r,��=AQ���c9	5���ܝw]���'�GK�� �e�(�U?�م�Wb������hl���Vu�HT=eq<@b%�w�ym)�����f&/�၌D@��G1�m�<=O��@��!�r"ն�VAKinL��ƞ��X4���'��䵢����lQ�;���5~��q�{�1TL���፰	����	h�()h�ʝ�?���[� �����ڮ2�v�|�����hξ���O� f��w}��q��	R����l�
�/]y�7[h�g��$8e}���(<XUʲ�CQek����G��Zs>�jԥ=f��3��&7�0��H�{cUv�����;Ñ�ܰ����%�*���P�������~�L{L-Ƒ�Z�d�������z��S�YxԼ��!��헤�[��hC��4�x��v�\wS}Z1�"ȅ�y���!�cbq̇���(@jqT$�G�ՕZ��ǙE���5�hoXN~wyR1\���W�i��\��@M��������BgfV%H�l�礲T���P����#oSڳ����
)����&+�+������������L�ǱxU�����i�������%{S����g�\*�()�΀м��]�';|���"AY6�O���Ch����d$f�.�yj3T��/X� ��>>��$J�X�l����X�+,E[������M"~�irg�$1�Y{=.�J�Ȕ�~c�iZ��w\� �E�)Q��E�WBW^�,� 4doj�d��}ÆNt`��Q�Cͽ�z�I��=Kd(�R��0'*�:%��b�#ؿ��\D�1�ZM�F�Fm>������O��|�H;V��h��;L~E��L ���V;fn�<I�.�� ��M4��H�2 b �ٴ��a\V�B2����Y�xh���%�0���'f�~�Te��G���5���{�!w�oCW�Mt�ț���"���n������A���S�vfI>A�_
��b�i������K�K�����1�c���Uq��AO,�����e��w�c�;N��Ӷk�6f]���B��M/`iD1�D�T�?�EЅ��LpD����:yq��m�H��{�4;��"W^�,4��L7���0��	��,��-�� �wާ�r5's��0�g�;���̈�
ʀ�7V£�#䇾B]P���Ο�Ni�a����Ѩ�:lr]﹎Y<��M�m�Uc:�@��h��<Ih%gm*<]�<��R6�E��@�S��:1=����ίɢ�	��/�;_���Yl�nl��,&���䜕�.�oW����}��@���M�]�j�ߎB�#e�����2i��)�g�Zr�i��]^zb(�}��T����Td�L^i� ���և����/A&�����1u+sK&]��#�O���K|ץ�R���b��E�T^͙_�x��k��YK'�yg����^p��Z !�|c�YW��" D�.g�dJ�)�=F��~u�=�F�MÆ���WAr���ɬO7����"�n� k�s���~ԆftM�*n�@S�i�]j>q�,ri���á���I��sH�����Q�2�u>W�4l�co��]��H�@��n�yPQ�/:�KS�[��o��_f���UO�u�s�����������2n���