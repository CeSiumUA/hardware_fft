��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�g`�vQ��0!mC _�e�� �ý�j�
(��6��N�����V��iv�y��a�2@����<�}*dw�4:Fd443���f�[����*��g�!�`f�ޚyP�/5L�6T]��4�*uj1�PS�Usm�_m�'A��kB��&�M��#�ʮ�az�|E��C��+퇦��@�N��s�7D�-�ür8�qɨ�'���_�� ��1�lѨ�,D�,���3�ƷXX�����!�K�hk��Սk���L)S�%���n�4�{���}����� _�k��B�Y�$s5��'(����w�Djf�G�DD����$~5�	 �J�o���7+�D9�>�}�.3)Nө�\�T��<4)��>:1!�t0;�8��`�Ă�[%��#A���h�)��S��t�@�+[�$*�ffc\pՂ�z�}u?9}�E���` ����0�f�U�:Xh�K-�7C��v���'ò���9��X��~��Gk0�� ��
���pO�dX 7e΂��(��-٫���δ�����|�����0��C�����D� �œ�ϥ�G/�,���E@q��d�ff����K����b
M=�`�����q�<��*3��z��UE�?Y���1�j���S=B,-�D����Q}�P9h���C��n�xN�DIC��j)Nn���1���������6��X���A���0wC᷃P3q�9���}UB_�C�>��^}��C��oj�9=��`�V����dT5&�TO�mګ����
���`u��z�b�������^X
�/ݽ�U變+՚G���t.A@�,��q��뇋bK)P%\�Q�uH�׏��jΗ��_��R��P��&{���ɨC�8Q �}��F����l:�E�=�Վ6��-��a�hj��T�pO��	�4���w��'�}0'ёVo�_pB6���c�ݿ�V¦f��[WQ)u�(t}�U�&2��B�tqw���k ~�3w�:�E@Q�9�n���1�T@M��4,��4�S_'��?��.H>8�fQK�Z�C�ݘ�����M�>�]Az���\xAn��wg�����6Q)�F6~�yr��R�����r���jڨ�oOJ�@�ӧ�`Ҋ|#�A����E�	<���*?;=2o.B@}۱`9{G!P4�;;���jΩ��j�{���W�0�4An�TY������h/�	x
�4 ���Z����o�,E3㔁�\�]b19����&/�^�N�$�Y�+���!�<�xt	\�9̵�J��s+��fC��z@)�g��.7��~߲���F�q�!CP�?�p��]*@�9˒�;�wh��:&�wB�r����*���{KāM&�V簣^���0����4�XH�B�C��pT�S�΂<�9 �<��j]�"�Y0�) w���#QS��q�Di`@ӾԻ"��JGF��U����qIw9�g��G2V�R�,*��8O���/fkhx��rB�&��b8�RՁh>a���єHS+�Di��Ͽ�_)�ٴ$�P<2b��7G��,��|?j�,�@.'�A-�J�E��0��G�p��Ő̮�w�B:��]A�e>"� o��ߍ��O�W�FWp��U]J�H��͡3j3՝�
�+�*�7a����'�y��E�t_讟>�����1�ŵ^	�
��N="K��P��4��Tt�b[��`�3���~�G�ݲ� ڤ�dܽu)GGA+���ߕ�Hxl�����)�B��J2Эv�p9���N1uk�NZ5
C��C@�ZC�M�����8R�C��qN����`ꋧ6�g_��t#���-.�J�3
�Z��'d���{TKQ��)]�b{���46���(�"'t���ACuZ�1��Q�yh�i˩b�+5s��@�G F��� '�Ϣ�)v�;�w`]����NIu;(�#��4��JO���̴�Qvc�Ԑۧa�����YD��r)�y ȓ��F9�����&�uB�B�b����M[�
J[�����M'a7�U��[��\$A��{�kqv9ۦ,����R�!��hy�h Nxc��Po`Mu�M�k�J�\z���3���9� �����e���s��������p��0����v�T��V�뱒��W-�ټv%탫3^��5�|J����N�$ ]^M|oY8`�
���M5?�
�|��N�]��:��a��=��O3�]�eN�T��tc�4 ��F�~l�$2Ջ�YO|�{'�{͜��=�b�tEdc���,�1MA;{�<��`Mu��r4x�%��#t���W2��}IS�ڗ�PR�Y��<����ȧm,O��s����c��{�O����d>.�n�ɷ-����3[����_�,\1��/����T����_ƛ�؊c��Ul�0X�c��-���M�>�R~��O��`t�*�V��<�������T�f#�xb��j.���3�M/�7�_6������?	mo���B���S� �,<JP�{��4*��_3de���@��+>K��*��}<��*qF���%=�hf������Xk
��2bj�/� +, ��;N��[y}O���\�y��ߩ���<.M0N-m(��;d0�q�j.��B�N��>��%�M����y2�t�Ȇ#��5�ϒR��-��m���E�J����<���K$c��]�:�Ɨ�@��Mu���ܴ�zE�=�w���[��>�Ϲ�)���	&���%�DF�K:��R�.�*bS�N,么��
 �)�R�5�P3�A�����k(�?�~�k4�߻�A!�)�������7Z/uȳ�}��(LA����[��M�忰bB� Α�\��Q��*�.�-�����҃ԯ�b�ٸ���<�q�.�|��IF���ߕ׆�Sy~7�֑О0xY�p��g�IrD�����JcղO��=�ṣ:�~�d�-3���y5�\��Zt�G�ћQ5㊠�Js���>���r�YyJ=z�[�f"�24����`��qQ)�_d���B)�Nvn�w�uy���u�Y+�2�����7�#(c:���l�5ܔF?{tPj���o8��L.��!ǼR��Ë��3F�>�H��-�����ŕ�r�i/��7vW�w��:��z�+�b5_�]a1
�͆U��w=L�-q��Z����=x����cDU@�C�đ�״�MQ��T�@G�}t�V�J>yT�j>ة���ip���6/�#�f�,�_�t+O�)���W..D�E�N�nw�����(�6g^����YO�f�tjE`�ݗ�pSb���vC��vl���v�hO�ĸ W>�W)���_Ԅ���x�X�! �&���N�}���P�WY�N�P�Ta��FO;~�����q@�_:P:'��rc�J@~^M|@�T(��Y
X������mo��h��ָh����\e>���"B�EA���߈PV7ԷG���|�:ƾnO�Xr�Cv�;?�����D��YF%����⽀y�S�}a�����Veʿ�� �}N�o��?��NgR\&��=p�li � ���J�C��N���?���ӑ�ݶ��`�����a\+�W7.=Gq!�AR
���l:�8O�,=3��d6����v/#����� sz��*�Y�w�m���<y��9��� �{ݪ4���dz	���O��V��rc�gsԉB+TYT�Kh �
$&%��.�b 7��5?����kC��<\r�,\�R)/�4�u�ir�@MT6'q��S�_u�e?T6�=��M�K�Yۃ��c�w/IE��ޫ:�e�A#�^�W_�������z~��g*�����)�Y4丮��g��9/1�r��6@����jd�� ���AE΂�N޴N���'�A���X~1O�!Rx�9$���ʑ�Ժ?���~ΆFPZ�;(��2�S�k�ɉ�������\>���<�%߆*w�/9���W��E������&Y��yi�y�)����}Y�(��rYYE�
��d͞���;:��'���Ӫ��B��J��57y��nx�zvu<�HT2jFg 'H���J�����}1<P��4ğ)!�^�Ķ�D�U�yT@��DI�W*�B��ygI6��;l+�q���	�O��m̉��zS���U�S�dgb�������	��9�-�Nl�����vc3��C��G�XB �hB��^k���`o�`aI�S�'ac@Q���[]�/12tc��6e�K��D೗6n����Ѐ7�l/=(����ϱ�|���RuȄ��V&~gS�L��rg�G��V�	�^nK��w��M��Kn���.3������|�#}q�*V�NWkyB�"-�_�z�"�R�}���-*��/��;G �Qm�aB@ ��fnyo1�0�(��RMk��ʏ�j OU1Xa�x4�<a�>��Λ�x��R
��R��j �~�����ֶ��Wl}bq��3%�w�n^?���Iz5]/s(}a$Ϲ�/�͉��2�2��h��m|x'�K/V�k[��"���S\8+"Ck���u�> �Yp�C��fA*�"���t�?��
�(�M�
��LT���M
�i�G�P��0�M�˻5?0�Z� ��=�{�t_G���ج=��;�&K��k�����2�	���l��z����YNQ;�����|�z�w�':6�X�h!r�o�F)��I��	����O&�3J��7a���L��FV��MM��M	ܓ�e�)E,^2���Q�X�#�)�0z�G�_�DdD���n��0BP��#*��6������U�{��# �,�C��A�uM��e�d�6v���-�V��Ҹ��S���&HԿ�1Iϐ�@ ������}�Rv�ˡ���%a���VS$L�Zz���{S�]H=�r�P������Zܝ'/���wC&�{#��� R;���H�7�ã�:�2<3�^�\6��d�95.�Z<u�5y: &D����o�;[F .F�ِo�,`����A�b1�׃`�}�	�}��-�z����P���)y�0>z��bA���6�-/� ��I��
߰�_��h�^�E-�"���.��ߎ�Ka�b������$��#Q���}�r������u )1��SV�� (D���5�2�X���T�,��W[��dĈ/�&e|<�W�hJlX�$���^�y
��S���~m�V���:K�bb�9�:B�����_5�a�dF����ک1��כ�=�e��(.Sۚ����t�GUm�G7���|y���,�l�d�U��M���J��������zЭ�]��:��3B	}��VA��C\؅F���$��G�*F���RQ���?}Ɣ~��A�� ���1�g����ƞ�N�r�Va�YJV����j5P`�t�Q�Y��81rj ��]��p9of?��/C�}��u�T�.����CM���w!,BM6�\���&eaS�"�oc\A�r�	��,�WCH*���L���, ��:J�Y^�%c�Jk�w(��H�K����#~���Ek�ABbn����C���sy�ٻ�aO�2��8�z�����}�VI7oa�|˽T\��՛��
q�S9������.���K�t�*�gf�K���9ep�s���O�����L���`zU~$
̓XɎ�o�T#��3b� ^�ȦŮ���KՎ���s�6/q$U��y�H�/�)}�Z� ��׮�U�k�}�� GN)�=������z�C ����4W� �q�1��@J�S�O��=�+d�O黪�%L h�̤Xa�Lx�70\����b]n��1�����A��3~�+N�7����G蘱�wg�%0Z��	i�pt4��Ïv�fU�Vh��|�w��=�3�ï�����T7�CUx��4��KR�~�6�ȵ�E3�+i��&߱��|���kYe�'�)�ė�R�������̫�m������p�UP{88uM@��d���Y�������+!7֛��_�O�93���k�E���=bA�am_�
]NJ��A����@��}�X� �l�sI�����/���N���v��'xQ�O�� ��d��l�_�C66Z��5�뱩��z7���usr��iSY��Hk��'���O��d��7@R��)���(�P���?��<�H�6K�D�*���ց���Q�l��H9%��տ��x�r�G���O��b�����9��mHY�Cb-�Br\�ߡ*�&b�G��L���'CW(�۴�N�vϸ�*-�ر�7�/�-���_U�#n���B�~A�,�hغ��i�Ё���<y�R,�E�:#<U���y�V�MN�ŀ��7�B<���.��f1�@j��J�&�͸�t߯t�����:'y�q#��E;V!h�c�?r+�Xg�-y���[�4�i��Ɯ*�_h�U�w`_sO��u����{���-���ԅ;�ͳ|���C�_$��N���P�Q�tx�v�_�C�����9��]�s�E^[�>Y�p	��dRgh��߱��Q,4a��;��^
]�#���>J&~��Q${�jdgr�������B�j��F8K��)�E�I��;��n��]CQ��ҵ�/��H��1"Dp"�\r�����lx�.�9I�5�G�b��ͩ�u|��ґ�����_2"�ι$�^l�dїA�bp�QH����d�����i�1��(�ʥ��/%Ȉ�ʺ��3ߺsTk�
9��ʻwK^t=�Ј�dV����3Hvg�(�\	�<p؟+�l9�y*���&�R��ʅ��"5�)���X�����X?�!o�i���CGn=�D��8���N���)��DF��\���_pD��Y��J6�<��`��"�@L�?�@�oC��%�J!-�$�x�������0�<�*�:�V+���T�C�p8�i�c#�E<y��m�9|��p�������	���%��ݥ!	|(�����ʤo�Ё�-�c�q*ߎ���[W�,K"�����m`���E�@<���o�"cE:�^jUί��Ypi�%lzP@v��"��&c��:�a�Ť;yV� g�
	�t�$��I���?�'�1�4f��b�v�k�t�������K��9H�[���w�*X��uJ7+�o��_�Zڠ~X��`� 8�xUDǅ���vH�X=e����/�8Y�����)��b�~f�����_-���'�E͚�]Y����Hw,:��$onY��'&u+�+ޱ4s#!;)�Ƌ�C�2�-�)�@#/[��җ������Bo4��6w��!������S=Ou�!�� 8��ץﶾ��j�i�$);���Mi��x	kOu�*��*i�(�k]i.K�QY�� e��d<@#��殹`���υc�g������/[�؍��sw��b�8�n�\�II��&g|�!2��&M�z/-I�m�s�O����#򕾕�|��閠�f�i�]Ǣ�ΧBwK�@��?�&}��9�ѧi;�ng�A��\���ӿ�*&��\-�֕ˮ�I��i����o���� �{|�A����3p�|�mry�YɜQ��So<���X��}P+��7�,�!�k���(��y�X4b�-:)�8�t������1瘳W}NO���*�2hr)�r�ь0�.mxO�-9w��̧W�+Pr�1�ȆMv"�t�����c�I�#����h��3�������C]�e(��R�Q�Y��q���HyU&�)���U,nIm����P�$^MeX�i"���/��q�P�K��یO�	��H�>��n��|��̵t⑒����B�}�2C����������͜+��#ZP����$���3r�%�R����e��Q�c ����L�d7�����z���c3���=,��&���ɢŞ_��k�|�9a�Lb�b����o�a�%l2h�x�F���.x�ɬ,� ���Qc��?��z�Rn���d���tM q}=R�����fZ��v	C��JG�O`�ܶ	nE5B�����CM�ה����^�����_}/C�P�=E4�7���D��ia�H"#��;���sa�`���?�Y �m�-�;1���;����ӓ*� ��s	J��iV�'��=*˝��!��M�r#��x��� ��z��@e�9���k����&g�3U��D��~%Ng}7������n��@%��}�
�b
=���ۉvBF�t�����R/�c��wk�Z<�����5�s��B.{��Ʊa�p.+)�&˱�����k��1����>����uA��W����u����O�.��![��x��wӭ/��cLD����e��k���F��GKK��O��?��]��{�*璽K<1��>��h&֪��F�ۑuuo:֔��aDY�jϣ��Ñh��>�4q��Ă2F�O�7-�5$mf3��YKi7�P�%��1�x g��s砡H`�%L���<���mY�gƌ/�Rf�ONB�͚:7Q��<c��HO~��	��B��k.�����J�\��L#�;ߓH>�z}��x�j$�O$2Y�gI%�\W������(�C�����Q�0��>���]�5$��ˍ��IY���9ss�G3]�N��R�8���x� Z�a}�CВ2�kC"\w�w�%3����#u
B(�����%L��9'�.�W�C1�Ǹ���~�3�iA��X�u4��Q1���GjR%�c�V�sk��$e�t?���0���d@�O�cc�7��1���'cJJcy�!\���1�@�i&�0<?�Y�õ+3���Gϯi_����Ǧm4zЙg!��?IX1$=ە�->�_m��ܫ���@۾�S�f",: ��H�����2�y�B�%��v�><m�ZQ^�2nйT�T�fYO�S3������I�85�ӷ�W�DM_ĵC��85z�&&3���CJ�#zV4#�e��/�b^��������(�hݵ��ݼ�U�^	g|�� <[~@����\�Q�J���p����Q�'�q���r.Ph��c�ݱ�w�� c�W)�@UcW��S�$]�O�� �т$ʠh�e��T�:B�D`;'JkK��Z�C"����~���.���ܦ܄��x#Ăr����`7�T]?�+7���4�M�!0:��
7�K3���^M���f.��O���Gn�<k�yW!�?*=k�H!��iK}W`>f�@��%����%.����F����,|��s��Ƿ���6<!���Oˎa��t���K��T#�a�}��'O3ebL��{�O����z4IF����\�Q�,%$L ^^VvY9t�f��J࣑T�fɝO�oŦ�qX�$��΅����!�iO�����2���b[)�򻔌
�˘�5[�k��PU����2d����_�*� -�Q+�:��B��*�R+ ��&N �j}*����������p
�<~ߩ'��7�e��뚛� Kws,�v���X �,3���B��2�&���YЁ�#�gO�͡�2���8�f���	b��K>�o�����0�\Z��7S"7��.��i}�}���(�,��_����!������U�|�n�Qx{�?WgG�%s�ƫc/T��o[�nv��ƪ��(�u��fq+)�ٺ۲ڨ.㩀ΰ����͝n��U���V��ݸ�����ԩ��}��d��dZ�(�,턙.?<`1겐��c�8^>��J]�Qi�a/!���p���gD|��Oԕ^�VgXӶN���MB�*ұ�}�M��٪0�3��d[!� WLX<m�3�ڥ�sI6ϣZ=�.h�bz�1o��}�����5M�0�C�Rbw3w�5Z�M��K����_��ӓN2����Kx��k88�]Hl�h5t7=[#"�_�2i����y���m��
9��0u�̘����X�����B�ָ�J�@?��yk��ֶ���i9(n��}EO�/{ʬ�MFˣ�Z�׎<`�]P�ˀ�g�F~hۢ���3������m9ꡗ������˖Yd��n����������N�1;�x��y���̴��)��7l�ĵ�����(���&��ZUSEL����Ŝ�ƿ�sW�Q�5��-Fjө�x��S�nB�j�&���ڻ�!��㭄f�'�s�g��R��
�YC3+Eĝ;�V�n��o��庎n:�28{)�)��xJ�`�M������<�k�5�@�o����;&S����M�n�7A~Ķ���v�*"$1��"�q^Ʋ0��q��� x3G�̙�W�ua��~�}!���`O��I�}��\�����u5i��������c���M�� �x�=nI`4��[�;{�)����|䥭S�B�9d��I2،����ď��ds}������Fp�e^!���\��!f��of;V�+�;lE����/�n��2@�!e AS��u�@���+[�?]����y��"��W��֛�vEIw�h�b�f(��\g���(�Ac��Bp��ڦū���TF��u�&n�|��<1*G�2-�
sgP,��{�_�iz�E��ύ�ZA��u)䉧f8!���>�?��(�ut���Q��y�0dl���P�t�d��Z��Ir�Z^�<�)ֺ�U���k�>[Ύ��PZ�XJ� !r0,�78x����4�&�Fof�iu^�wjށ"��;G7"k��G��LW������&�P!O�G�)H�)��?@��ƒT#{1��;�!���t�:7��,��X�e w�J1r���Md�q]	�?;���n���)iv���ԟlRg�Ej*�)|ɽ�c,27���T<�A�S��.=o�^�m$�,��̐ɇ� #N���s�7]TM\��(�� ����D�y�Pm�fř��� 9�@�(���x�э��Z��z��������6c����Vu��"d}D��p ޭ$��ڹ��L�,wvp`t�<�>��P~k^�H��YrQ��	�K]�7��ɺI!����hz��rZ��!�41|0�t��+������t4�u�R)�������#[���I� ?4P�n䛮=rZ�� �_�`p����0g:o�g�d�.�b�@���Ћ�-�S�%_���,j%6��G� ��uud~ �rCY�?������,/��z~Y ��d��'��e&(�̾�kBiͣ<��*������~4{9x�d+'w�%,�gi�ZU����JfF�f�Sj�M7^4Z�r�՚�5�1��ɏg�if�?*wq�:��K��I-�����<��B0�1Ut�����ؐi3�rqu�1[�ǐ�rZ7�><9⅃�H�M��عY�:	"����o�7��L=P��M��ya�t]0���x\e��;�,����v)���6ǁ!�UD�	�u)@���<����Z"�*�iQ	���D�ہ�ns��V�P�(�	�;/��CǎV���ZN	��Z���"_��3�N,"o���Eŋ�1�'`���7z�����`i.�}�Y0ǳf0L�����;����b�5Vh�������W/�`t�~��5�(�n�EΏ�F����%Ne8��A`����0hDfwtT&��0��V�Kɽ�Į�6c}��ր:�l���L������6����rU]=ah|��R�d������
�<����)��e�9�8Τ���i^; K��{댑���������2;��Cl��z.�u�������
�F��Mޡ\��ɩ��BUޭ�AeX�����1���F������+��Ɨ_[�rW|����CAcXޭ��8�� �/%	>�i�M�3Ձ�㇩k;�j[�[��W
iB8u ~�x�DN���N�Q�]V�f�-@C���8����ۏ�x<��FE�C���>�?��z��_�`��{p'И�{Uz(ڄ.	����*������4z 5�k.=7,�fj�>8;EŻ����` a���pC���gW���F�1���-�Q��[��|]/�:�!��Uq�"c��m�j�hl�6.m���9�i#q�7g�B	��+�2җ4�Y�K�U*���,e���.5�bc=>Lf@���F~�疣�J$AX��dx�#$��`rd�2-Z�ـG����b�c�������"y��iD�g�@��#K���,og�@����=�/@�:^Z0q�b���aa�X�D��ȌsS�}�*��\�����!���)I�fj���v�>��+�%i��*��^�~q8���=Ӂ�t��؇��!��u�Nh&���)���klO�e�4	��YP�x���@�{	�I�ԗ�W�VU"O�MFS|�P';	��ڇ�Z�\n�
z;�"0�q6S��4!#�ur.Td�}���ڤ[J���GIy(Jy�-;���R���e2o���9�jK?�qO�Ma�C^%���F<3��eؾD�<��V�:� *����Ύ�^�JZ���dM���<���l�7 �aM˄��j�1	0���'�ՖX�F�W@�8�&�	o���d�x��T��xȑ˰P#}б���\�7�Uw9�Osv17ӊײ�X��;���OEUQ���yD捞uB�pVf��ļ�@W�n�4��°)i������ئX�Q!N�=������z[TK韚��=�s@N��N����>���&,�>�("�S?P�XZ��ag�Tp!$�l���}1�Ň1�� �˱XG�,�#�b��Ş6d�f�Z��w{7X���Y��i"v%�5ߓ�f^��:�v�f8u�Ϸ@p�/�٧>o���h��j�2��0n�fS�=o�{��9��wX�?���G�T8JTk����q�`��#��؝��mSO�g,qh*�K�|��(C�狾T:��oe�^ޯ��+^�՛���;Щ� ��Q������"N/f��\�߈`"�2L����Gb���N+f��� ��I�?i�����𲺨�W{�܃��4�q�i0,W���}���U� �i��BN�V4p�0=���ų�Qg�d˼g��O�`7B��ck���x|fG��pl���W�Y	�+�(�;��?*z�G��<\
���6��q�j���(��L�(�>�6������Ho����i��N_YHW�� i`��T��Ԇ���&"��S=[����F
��y4���(t�΋J�{�]�}_l�3�[�
~���^U��X|jc�jn|��ǫgI:��X�^ � K%ƌR\m����k���s�q_���Y�K��!�q�Z��?6�^�a}}�Xޟ�������K@ {�"�cԕ��<�9ku�pu}"M�dҊ8�C����#9U�zwK��	����p_~��(�+��S6��c�+�n[�n��y#蒕����jg�D+h�ռ[(؝�Nà���&�,�sTQ�=�>�朑�"O�+��
 qF8ԓD`�y�-�]��0����m�}_�]���|(:���qH�\�	��⺡�i�cľ%�7L!��]�S����#��Rp�ō�*��@��/7M����@k�
 $V;J�� 2��N�B3��b���}��q�|cF�BM�b��vn�5Ech��bl7l�Ι��׋�ֳUʛ嚦"0p�T��j2��?��Ǌ�f������)1��N<!"xl��z	� ��$o0Vl~wj��Шv[&D}�dA����_�:z����'u]�����yh����]�(�MZ�f�m{*ʗ�+�{1˄
�C��A[in{:l{/���-�*O������s��U���OC���/UIEw�֚q�v�'�<*�����?:*3���려R��=�����\ �t(8x0���l�kƐ팳 ),�g����i�Љ�Q�7]�q��f�pZ�@�F������$w3�f Tj�A���!kVm���lI'9kÀ ��F?ޔ堇���pm���q�|���k�L4̺��_'r�ے�'�pP'�<�Q3/�麉��زODZ���N����L9��Z�ڪ�.�A��`�'T ?ɰ���@���a���7�(� �(��H����em��tG���:0�+_��OI��Ѓ�q	!�A"䵘�OD=[Z�L���K�đ�� ��*���u�m����T�i�l�J;�[���>�����f�%�˺a>�qy�|��� �جbPD��'�e� a �5�=Ά����;�rpw�b,���2�����5��*���D�7��_LJ��*�2�פ�S̒���]�mͪQD�9H]r�﷬�#�KR�n�izԇU��7���`��K~[���j:�?U̻-2�����c(��4	��<�?�Vxb�c�ʡ�d1�"��`�b�n�csE���� �46�Q�2(�.>x ��ؑ�|j2����&�� ��6C4(���筩�)���~Q	���F�V��c�j�f�%�Ò�;V���eN�@D����_�u��A�"�#�dģ(�O6:�mk;Hۉ�}A��/J"&uT�4�c�K�wA�����w��6���7��c�u�x�(1�Z;�}W2�Q��~a͎^O�T�{l�����%i��Av�z,V-��W���S�R��G/2{�. $�3���쮕7IyS�q��*ߨx�2��bM&�
��Ve�S�w6:��~�����v��ۛ��E�B{��HvM[����u�ٔ��׮�N��C��Q�Z�X1ZӡG"�?�hleK|/Y?`1���0d�E�!�I�|��"�?؝{��1yRR@Jp�xY�*I����g�о��{5-|����k�y�p�_s^��W+����*a>��\~����.��ʪ���,`�o�U�uDi!p�/=�:��x"��
��wU]To�m9�B�;j���>�F��%� �qe��8��u�"�e@�6[v:&?�[�v��W�%t���!��A��g6Z�&z��~�|
7����z���Z�`1�n�k���,)5N��M�L���kt湥�۲YZ�CGvk_�"���=�0�Ă�=�����*G�LW�6w*��*�j�θ�u�h-��*��x�o���4E�|��x�p4Uu�.D�h �29>�[�Fm�나�����K�\�γ���_���s2~�[���)Ǹ�ې?_�ն���.��b������_9׽���6�M��~��of��ŵ�&�q٫0��ȄZ�W���(2Ws�gW�>�^�{M�KCt�W�M8�
�q=I��Ej��\�ɭX����ݮ���@�h���(<ᵠV'c�?s�}D�h8����
�)Т�iVrEr��
3>����C5.ˬ(�'!��lpFL�e��ӫ�A���Y�3�C�~��Oa5��"�ʪ��nL�rdW2�P�����Y���Z��WLK,�"�!�wI7� �g�I04�,���WNO��.o�F���2��÷�z�ö��f��ª� �ie����l����g-�I��8s�fiN�Aġ�]�/��`������s�k����g���V�|{�``K�ݵqb�_��z@���k��&�.��;E;y3�Y�������Ԏ:L.ڠ ��,�@�_��&(9���W��vQ+�Z��t���D"�w��a��r�Z��B���*-�)F�B�2иw�Њ�^22A, ��yX�2�dQ������� � ��r%u��K�)j,�l�2@�OhK���d6���㾱?;���3R3[�{�4������#
��]N5N
���� ��MCfz�������ȅ~�<`!$��`��i[ˁg��U/){(�N%:Q�1㝿Rv �pA���6���-ن�)[F�`�բ����ϔ!}����{+�w�Jz�u��Qw�1��A_o�Ly�5G��6�Ҡf�o1Ci#�# ��*�7ݳ�VJ�b+|W���wؓ��`Ƣޢ��+�]$ь���k/�M �`��4^m���~���d3Os�*�R)����OKi4�b)	���	8�'Mi��RM_M/�F���gކ�~k;����$�����l:��P�Hji�G�hUy��,�����"����x{D%f��?Hnw�/K��'���	K� ���#j����JM�����0�ˬ��Bi�~z���h3N����;���Jo����R_D�)q"��硜�e&�	�u��	&�\����\h��(I�,d�W���v>y1��>]P�Ye^�Dyw���o����U�?�0rs�[Ω�gG�S�l�iZ���.���\'������-�W&"�i\�h(N$3G�*��Y��Ҽ��%wVՑ���[����QE
�<Ϝ%o�Ϲ���H���7�w�Nu��3����	�6�����l}52кm�fI��4�Z���;���(�,Aoqփ�ک78�H=���/�Q�J��� ��Kl*�y\�?���I�@[Qk����W� ��?3�:ܫ��uo��X%��V�Z7��p�6�L�$��������~7�K�,)�$r�ן�Łj�Q��Pc�้]V�n�bY��?^9} �~�<mOt �dO��`\^Uz*��-�$8���:f��L׼��i��j����|�?/֟g�n�m�����&2fz�c�2����Y�4�����\i$�$ �����Y���|L���g�x;�r�^������xuk�2cOP͏K��]�J@J����SZ8��T����3�?���ؕ�e}�E��� /ˑ��������v��'!�W��aq��ި�͊=�PT�����3Qn���5�'4�rP�#V�����i����#�-�N�'o�e�[�t;�$�pU#���{}��!)f��ok���m���>\�a(��U�As����,�<�ˇ��<���M}�^��
倒H���+�Zr�����O����b~:���Z��E��Ի�[?�GTi�d�q�������LRaF!jV�4M��t���ҟ��	�q7*��|+~�갓կ$���+L^��Q��wҎvx�����/�ɣ��},yǂr'���i�Y6j�/�;IR����e�Ņ��_�&A�M� �������0E�d�r^e��������HK�Na�;P�`�ȇ�Ԝ��M3WƔ�ʇ�W{p���K�2����m$��r���ɔ%�?H�rK-����^�5�H
�E�1�����k����Id��5q�~RE��D�ɓרTq�\Rk�P�V�3�gّ'1������a�rD�&��G�.Ss����eY�<�UW��h�k��,�2�-�����uѐu�z_�,g�
��p�y'�8?�u�Ȯx���c���Y�p�%�8�B�>R]�<D��5���y�)+���_8H�8~�a���.D�bD����ۑ���zSЯ����z�S�,m�,l�^K� ��]�.n㄃���"���ԯ�'���,���rJ�q�V�B#���E�+)��KgҺ;y�G�b��q-=� � x�+Hm�����`����z;�ڂ�����ЃH���V�E|�OD�]�.d�ǜ�ŮI�����f3�n}�n���|�O�vn����F�E�tӡ>�p��J�M	��MkU.��rl��Q_8i�aA�D�=G��V�O�H�n�ZXB�*V6_����_P�� be��1﹈�m����ڹ����$T�.ޚ�Z9��c2z |6�`/��m�3������C�U��{c����~ӏ�!�rj/���5�O��J�M���@�r��Dߗ����WE2������L2}Ry�����_\��T�<�})�p/��a�l4����&�Ӛ[�(�Q������DYS�w�u���Pϼ˟�u�߿����3����������>LrV/�{��&S����Ȗ�\B�2M���_�-�WZA�w���r%�S��[6�V�0Iu�b�gJDeQ��F_lu�֞q�Q�������L�/���#��K��Tv�X!�o%�_P[�d��k��QQW�Yݴ�P��m���x�w���~�c8P��$I�B ?��<Ϯ	>�K�n�4�1Sa���L[�$%���k]��%�?����S���=�{��o��2y�6B��fK"�zt�׃#}m�#��״��ۼ����'Ĳ!�J�[�U��T��K:N4�UH�ݦ�z��@f�{�9o�[|䘗���ՠ�3@����\:#?�`䓙㰽�z��5�a��?fЪ_ʪ-A �%u��r��1v�����!i÷6��^�6���Xk�q��P#	)��?ۡ�'4a��0zUv��Jff��=6����ۑmxҧ�AыA@�RmL\�T�V�!N%'P&����V�H�ۥ��@Tp؃<���8201=~���J4R�ل�X���7z�?�XJ5���R�k�*�P$#�u鈦��(Wٴw]2�I�dk�ԩsmw	U��b��V����-����;{��>��'!��s�ϐ趤��v�F�G���1��тտ�&��]�s���C�|]?�(�����E�\Jw�d]
B�-���R���)�J�ZK��:g�+��]�����N��׸]�K�*��S������0j�HHhzH�`4��qpg�W�a���!U�g��G�8,��BH�p݋���ֹ�-y��4RC?G�'�e?��V���o��ȉl���n6Q*	�/ST�p[۠/�b�y�]���A�"��f�б���;R2��'��&���<�&Ki0�5��@�_���j�����Ԡ�_���.u�W���Nh��d
�Q���FS.^T�۽�DWF�u�U�9������Ս��W��@;6Ӱ���.X6![&(3�\��C��=�����Z�"GG%B�-s�H�uY9���e�H�/<�]k&Ҏ▶�?u�(f���em:+� #�X؜��ڭ�Z�r�h���g6_��E�d�kTf��0�F�Ny���_����9�b}����
歑)�5QqB�b�Z����|aX�L��H��"5-H�{ ϛ�Q�tP�n�	Z� ���!UE��J1����{ ��8�w!�}�����:�֩=����j�(V41q+c��m��9���˥��p#PPjf�=q~6�01o"�E�2�=�w]߯� �썥mFLqo���Q��˪�a��66�� '(u��(��#��,�A�=C�����x������0���ɏ��HČڂ`�7O�z�7t��'�)b���`��T3�����z�T�o��[+�R-���&1�y
'"���h\j9���'��]cKf�6��x{F3��9�� �b�B�g���V�ͷ�h5��5��s�F�����b Yʦ��]�Ē��t&�x?ӏ֌�ν����Z|�4�X>b�(G�N��K췕W�׺qe�|�u5�A�+�E���Bn�Q�h���<�K���3@�U_lK��.��_#B�Գ����FC7����a�쌕���Iq��# NF��T>���L� �>��^�m�|݉���4�y�m4�C�N�w���h-t������	�e̫��L���	ꕦ5U,��H�{:�h^�y��>��a;�^���)�>qL
n<�ѵ��Ѵr��j��p+�p*�L�A�k;�<:�����`�:�e�J�>�,�qSW�9����g?@Arv���i+YR��#-��Hр:߯�0�N��&]�o�X���m�F]�z�%�Bz�Mq��O���2�_O?��8:O��jC��?��{�����[����|s��L��	x'��@t��ΐ�p{&��"1��a�-n��!?O�g�6Op�i[�u '��a��z�t���V�_�GlC�Vq��F�� lLI�.����+�݁k�~�:�׬��B)��qD@f�A*F;�=��y
{�53��]�K�N�`�]�'0p�R궣v�-�� �.�j��ʤAYR^]{˟G���;9 Bҳ�Lb�(��Y:�#o��Qp��Yחg��H�������i��M�R�)Sƚe/K�b�*~����6rƮV�^�t�\��\8���er����L�}��*��ڼ*u� �A���w5�W�̜E����h��|7�)^�r���[N���b����J���Z%�{�zG*����js���4wj:˃�8��~IX�XAJ��gť%6ʪ-�Kc��w�#�"��l���e�FŇY���c`�h����낻,�q���?-a��Β#"@���fuU_���2�q}a��Js��ՍPu�V�B�&�o{��p\a�>�$K.�^�lM �z�֟��Y��A�#ꆦ7^�u�q5��݆d��@ݗ|ܒ���	��*饡Gj�|>��f#�� �p���og��*�}�iݒqD0\z��h�bFgq��>�u1]wXQ�*R��Dn)DY��Dk�C��Ѕ�QA�N��	����k_�`��[�ܠy%�U3(A���lpn�VU�q��`B4��ݩ�e���@��i�3s>����~x�]v)�����|�����Ǖ�X����.^Ĳ�+���O����O�[T����}Ec�S�D8��h�����/!m������ڍ�܀D$�*�I�i����{y߷���NZ¾�ύ�>��ϛ1�ڈ�Pt',���'��5��;{�B��ί��{�U�[Ј��4ITg��)����:�W�Ǚ;"�m��v2 ^��a�ޙ�P�jt�ɻ�dy�4��o����w����T���!�����nW߀�9N�%�,p�ǻ�X/`*Ӄ��7��0
�p1S��ɜ8w�_$��p1���C�B��o�lK���]�J��������l���xG\�:�V�=n/*��Y��൛�E�8�:+��迁�9�!�&��������A۱��Ֆ��Ci�����&����b"W�E��%�Q �Kx���ؤm���j7��=�>41����e����[|��<�1D�W`�M~4bU%��;�-�:ˁ5���f!S�
m$կXA�2.���y���HQ�K>p%'h����=��|;It���.��dKF�i�{/�EV��4��hM����n�KM��F��5������7��Q�@��Vt��f�\�n�Q�m����}�[o2s���G<�c�&v�b���/,���o�C@ �#e��b:߀�J���]����.|����C����]5�)aF�N����e~�,p9M��圶F�f�����P��듺k��X���X��Rxv����㗡S�5Q�bC�\Uo������F*0�gj-dQ-?2�QD���ܐ:�a`�p�Q<�un䓲ۘ�L!{�G.R�D�<��V'|�y1/<enn�9��Ly���0p^or�4��=��8�)�;�J�h�/1	�S��X��:ԇ�0!].&�l�/��x@#;��,Zq��_*ԁC�&�������������dE��Fg�}8���N������/s&V��4��E�`d]6'-�\Jwhx�4e�X쉛�X:�kxڃ����Z�e�cw��]M�t4��MÑ%������3eK��׋n��<����C�?��r�� ���v�3* Q��H��p�'����_9w�U�>�9���ip�kٿ�Rr���*�l?�uD� aX�
�oԚil��\ط"�H��J2��|c���PR��;|Û��Ɖ�����ސ����\�/M�JRQYx�.��h!&���*�ȫ�vz11�c��l����vmi5�Y7>G�<Xה֗*�f"{-`CO����7%���3��wa^d�i��Dq��l�d��r�%
�T��"u�y���j����v��}��B���"9,�y7l��o���:������)x	�U���9��E^��y'��+i�8�)�°<hQaksǨ�Fܤo�-_˨/�*�̧��"�S<��L~B�y
e�+�57
�v����6W[p��D�~�_8C���~{�c�)���
<��e���?�\�-���}��{J���!��^��]��߄w�7Ak�?��qoOŊ-q��V�i||��m�0�����U����i���e:C�h�^Ն�dTF��w�`9�Vȩ��ؐ@u'�1�n�{rK�.(��%"4?���8�47>��_��~�|T�ԩ�W�=��K&��q4��1��z���.'��ז�#�����:l�?u�J�fjf9�����@w�c���X��7 Â̘BK�	y5Pi���/��w����ҡ���P)8��r*�� j�EҸ���:z�K�E�����2��K�3\V$i��ֺ̂����h��-'�挙�P��4`�èݠ�ˀ�������d�r�R��;�ځ��^��}�J��?�n��*B2T��n��ZM��"��8�ڔ"����U��ۏ]�i�Ụa-��X��c�Z�+�џ�cO��9��8b��j��J�_�Z��ª��c|�A=�����Э �VVn�#���!V����s�\H\*5Lec����g	i1����W����٦mq|�]2�D'}�\�g�KF��|ch�t����O骰=��,���x�!zr�O���*����e,�HAn�y�+W�����^T��7=r��Z���aT(2:��ԃe�~���o��X�m��!���;����˲��>�'�P�DMJL¶F?#���w%��!U���W�5R���OiE�}u��	P� �D@(�ZlZ�UL/�c@���a�Nb;�,���s�Rvv����&��ʭK��k }ڏ`��O��T,��{? �x=&�;��[6gtB�- /�x�ۭuW#{��)���ɤ3	t��E�-s��^'uF�����@�~af]\��Lhx���Pͫ�����yd�I�*�ÅϞ�������W�ӄ׿2$�Ċr�� }�{L;�m0\���Տ�p4B[x��Z8Q1s����S"��z{&~�]�M��V���N�qq�f��H-)����\��6V�&=~q2v4*yi�Ĝ�)����lɪ�~
g!�[����L�H2�&��د�����0� o1��ry�p�̫��j�'�n�TfmZ���'^�K�2`��:�cQ�N��Ng��6�=�w��E������}�:�_���˭�h�!R��Vr��G�ҝ��Y�Z���veA�	��A��Դqe�2�޸��u�w�"<oA�Y1�d�zB5eXU[�d�0��H;dTpuvyo���$��L ���@ ���s�o�)'4�ב�D3L��,�KM����}�ቾ��J{����co�=��.�]*�>��h��GPԄo�����̟f�냅��VܮH��R��A5��
pe?�H7F�����i3r�������_DD���7;�S��ȭQ
��tБ� "2p�q��#ţ�7Х+f��* �{���G��-��o�1���AI/Dk�����3���̹,`��gP���[�]ߑ��J�[M&��z�3oa����/�C3�s�t�b�Y��`y��*��p���6o��>Z�s�k���([(��A��Y�S�Z/gh���'�ܪ 0��*8Ho������\�'�����b]��<��ۧ`�.DHW>܀+� p��<X��/H��Q���� ��P�����M:����.�%�76�W�������S*�h<@�Pg�n ��Jƌ�K�s�`�V6z�^J#ճ�=hB�hfa��y�z���bv&S70�8z�����������W�
���K�:�Xr��
K�@.�Q	���\�e��m� �O`�ȵ����fzǽd��:��4�����x1`DHX�u��=�����׌���6���t�	
������'P ��}]��������mj��C����Wyo,D^�����h�ټ���J<F���[��a��R�����b�n%�n�z�%xJ�I:#}�ij���=��|t���t��(V�V��Ls��U�������p5����l�����ނq����(7���_zM?�O�H��Vq�y� ?��t���5*{M��5�2�Dw��3n7پ���h����h�C�H�uPID���a~  �xZ�'>qk��?�V�����od��谻`]c�W�8��:���cHe�{��7��Mק��yx3Q�0�ARo%A��M�mC N�;|/�����e�r��%���&c7���d	��"#�I� �b�b+��޷o�����QD�"�=%���"�/U�=�dnU�6�R^�8<�ώn!��Vdr�����<G�?�����)��"=�Rs�Wp�R/��������p���`{�.rY;��l��C�ca��PF�E����N[��m#��{3�\�e,u� r�]��f�ܭT�p'GvP�@��6��Bڼڢ�]/���Z"@%��0�[ڮ�����|�P��
�}��Wo�r�9�6��T�*iP���|��?�3l�@dJ_ �����{7 �qS8��[2�r4�Rp����N�N��5_�	>'���w�(��p�rC0�&B���k]�Ʉ�o����@�׭�-(��";����O�H���W�K&qv�b�G`���{6���'�$�5�l��$+�dЦ��-�=�:�z- b�����O[Z�nQ��n�k�x�òy����'�|�J�"q������"H�p�D�+�?�:n���-�<}	7�*^h�X&ƺ��+�s���� zΝ��v*���1 �b��{���$�&�QI��m1�K:��B��_�i!׏�*d6@�kp<�Ya�s������5*P8;lK�8�~v��e�u���]V�r���$0��1�f41� �T U=f�I׉`��{$�<J�KG�W+��Ѥ��A��	���B�#fq���3�h�u��	�@�Ѥ�'8��.��tf�EZ���sY�����
��yL5f��.'�2��b���������E�žv00:đ�ѱ;�סּ�R��u<o�r��^g(T��Y�IB��
`S�~��
q8:ߍ����HX(kT;x�l4=�#=U�UmK}���]����+c���h�N`V޷γ�J��u�w�،�*�ul~FMY�zQ�;��7UM���Q�>��kv=�Q�BN�	,P��95k��_8���n�y�K���B�k�%ӝ���uϛ5pMN�F�ǵ�&�Β��$*}v����a��}|2�ׁy��@3]tӪ?t�p�?�'�t�F]T��ˎF�$-���	�!���@��{dD��k�&\g�K��0o���8��o4W�����.U��q��eI��HL0��3{�U8A�(V7b�c6_^:��m�x\]P��/Ъ�ƈ]|tfes[k.a���m��M�r׮���mՈ��$kV�mꢃ̷��]qM���ؚ*2���7�Y92G}Y��j�N���Om�5MJB�9��L��������\ϕ��:u!F[|�����K�&��w�Ə���Cۛ���O�<��3��\��g�w�LF�o7����p�6ޛ���x`�@�x�Ճ����d�?z$��i'��BF9�W������g�	�)o�P�r�B��?�3
lh8�۝`����Gj"}��p�Hp$g�u/��)����QE��W$i����9#�Ť����#g">y��\��"YMv�c��ȓ6m��T���!�ʙ��rf_�aכ*.C��87Iv�nU�D����}3�+�������}�r�)ў��)�RLQg�% O�%�VO��d�#�[k@��d��-Tm)PlJ���y[ꁬ^�Q�$����������gP��M��A��P�\R�uh��$�TA��d����>SJ�8�����w��j�"A fP��n,i :�k�^��=�� ��~ş*�D"��(���7}O��|�����g+9���H�����Y������1;z�H��ai{Ϛ��!C󤸲�^�\Ӕ%ܨ?��%�m6�^��y������n��	�Q8/�HE|��x܋�R=�+Ha^�L��neI�R�b�3��cvm<<��W�� ��^�л����(3�X��Ha'��L}��ň�N(�W,�T'��{b� �Og5N��R��� ���~j
��H�؃v3���;Sk��&��4U���ٙx�)nd9�t�2$e�G^���篜w��h��Y4�ԛR�V��ʵ-X�[�>Z�A�T���?��o��Uz z.����Cy��'����r�g�P#ri�Dbai�d쳆����������msH�.��%Ųy�t_2���L��qC}]d�*����*7G��|��wC��:Q�.�(�J���@`�
�8Z�%>�e�1��YB�$��3���k���P��Hph���P���ɂ���'e���ܜ�����'����Sz��Y��q���^?n�Sek�,���H�<�&8�"�l�;��ĘRLA��M�%��4����X9{`9�ڙE~j��z�v��3R 7�� ��?�9y3�Xr;��8����l�o���>U�y�|��y��웁wx�M�p�$9&�9�'��0���D��4�Mg�/��K5q��aI��aP�ܦ�V�q�Q�j��ɉd(x�շ�lU:��- 5����0^��\�h�-�%���`nQM2�M����w�-��j� ��57���>y���Hpwa�<|�2�\�<v� �(��2��ε_7>�AS�gڰc�ڰ�n�| 7��Z�a�rw���`U��O��#j���`��(�L���=�Wumޑ��c�of���I��s�T���#*V�|E�q܅>{���e��`M�ƟA��;�.�������<I�>�kY"����@��.7ܶ1|}t�I��RYI̫%�ʳ7�Z��l4�_jf51`���Z��2]Ƚ��]��A0�o@���;�	�6T�1B��M&x�?5�#%g����V�(#Ջ�H��@��5�v��T�ӵ{�h���n\y����*+�4��GaD�,����)?'�
��YY,����洈�xD?p��'+:�MP�p��8���.�#�5O���O����4�����\1�*;ڔ�D´'y�(0fG�,�����=T�8�eN#O
�o1ԫ6pf�:iȵ��	�  �-r�ȝƏ�DE�Ȗ������Ė�-!A�}s��O� ��a0&0�ժ)�����'kB.e{�d<�<J���
��Wg޸WKQx�D%�a��;�~��j�c�M�/c�O��\�:��e���R=����q��[����!@��Q��[x���l�J����U���EQ����H$z=^F�+<	����t9�bW�a���߱TR�ge+��jw���(��-e�0��1�-Z����3@�"�DВ�[�%s����^a�Dg��J�����Gn[n2� �D^D�ym��Q��e�נ�ݒM��Ī��E/�v��޽8��oLSe �7C�7��Q�z��Rk/B��� ��)����J��|�gW>��r����"3-%(=	�{���4�p�"rg�,�}ԋ�oi�,+���Kl��^��J�!P�3&��	u�a�����6�KD���:�#'z
��up�^�^؃SYm9���f'�?��Z��N����9�HJo)F�*���o��Rm1�_)��l����Z�Y�[�mHU��G&Ys'~gJ����M��q�%����܍�"�3+�e&R�Gj�T�����x�9�c�[V���y�齻�O���1%��Ǡz�{��s�A��:���+}ծ�yZ�9��9\S��Gݶ%�ζ`��(��"/?�����[eƊ\b�bQ�N�j_�	�%�	�T��p �������R�^v� 87��֝p*Q��Y�N�ޟ��2�vbb'~3x��R+�K����7Z�
@�\Vۮ��%&���oA��VD�~#�����ɇ�9�q�<�f���Oȇ	�dt�;�z㤍�1�N{-O�C$���̀�2S�)�E�t�E���܍�}@��bi*� ����������1ڜ�~B���̅�N�uM*�/����O�G\"���Z�4��
~��3k�%������}V
$0c�L:��M�a�u�K,�B�jF��?��5�yQm�B�
l�҇)W�"��u��)���~ړ�B��{�K0�,��S��:Ͳ��Ya�2F��m�����RNb�t�ʢeM}�ц�U�c��<a����^ ƚ�M�f)O:ͭ�&������3U����Ĵd*�(�?7J�d�h��`�{`gi}z�R������0��F(��T���G��(�:��n7��J>hc���5c�δ��ܐ� /$T�А R��<�4	��Q���g���tB�������@,�x�Gv��#툍����*Vv��e�D�g�ǆ%��u�u���Zh��x~�/�Է�O�-�?�M+5O��e턴�R�X��>�:�������N֧A��f"o
�d8K�ΫF���\"��)}qb,)Dm{@�FnD�])/��	��&"H���]��*+t��%|,U��L���/!zr/�];:U����5���d�Īz�/��s�Қ͂Gt�"���:�*��Dp$����+��&xq����pB ��퐺x�#u��Ɠ�qA,�r����ptU��w�t�QD K�$T~��E��lK�1��M	����FA�ʓ�i�?�C�_�;Ia;Aj�R*		��<����tr�J��kG�hڦȉl8��7ʽ�ov�-���*t�d�f���/Hڀ }�Cݖ":S�� ez�y- ��T�?4��6+rw,�<���Ph�4����w#��1���	Ě~�b��wN�NO�k�c|.H8��2߮�ɪ�K(g�2P�P�����S$f|=�S�������io������^HW �
��ŉ>��Ǝ�n�&�%��vd1�jQ��f(r�[;�Y����a@���z,����m%�m��˫?&�'@[ѻ�1lyj���Ȼ3*���}�zS��h�sL�NW�0��!:�{6��y��g{r҂/h���EL���2�r�ɤ��k�Q��ް�*�T�R�Ґ�8�-� ��Wd���r�O����.T�	���x�^s��o}�����u�]YD�9�n���A��:;���f�:�=s��N�/��
=���'�B?o�3�Q����j�~�u�-r_��Er(��Éd�P��t��pL�y�b��5����s�"{Ȧ���0U��]���p?G������4�����N��;4&, �A �\�S|�.����(��;(W��M�Ռ��N�W����a��V�?�lu8��bzV�+�fR�LQ;e���������_� �?��	co���f_������"BFp̯,guӎ�L�>X"]�R�[�ʅU�qI:���05R �pWU�\�<��s�}p�"��И�ҹ����/��jR�/�j<@$�w`[�(���qkPrs������ڮ��S��"A8� U�ù^{�`Q$����⩣.�+#��y��,��eKR��91Z�����(�ݽ��3�������
o��:@��)��/ok��T,DE�x��2k� e�� Y�	B��	�כ�k�@�G�_�A�N��q�l�S���w���r�dtU\�^k��k2LM����iD�l�����n��-a0wpO�
�.i��ұ���|?m�|*����8Fn_��� �6��ŏa^�]dA��p���'u�&��-�0���VwAw��q��o���� ��ϵwD(qJ�E	��9Fg�<��!�/˩�[β��f��$C�2NϘ-��}�=���yj��)���(쟐��5	�)�P�~��S��,�Bq{#� �N���3]�������_�ޜ �܅6��(4����1��8覽��w�:��f�k�\��<0����~ZJ�[�Q��<��	;8��܋�i�h�z�á��S��q�G�V�&��!�u�?9��N�8�Ҷ���9��Z�8�#���瓯����o����`�l/�P�ћ!	�
�f .����3i����M`u���j��,d+[n���@�s��A��/��ߺ�7��D�y������{��ϔ{����9�t���t�vn�F�+���t>G�����'�^��<zsBq��ȡfE��m^�
CH��J��Ҫ��1����G�+M�jq=g�c�����U+P/�gȘ\��c����ǎ+�̺nwF �f���Ɗ%���JTD�lF�'�����*�ժ?��g&�ghC ��/�iK���-�Zj���b�b�u�<|�eA��~�E���S��OSZ-�r���e�����1f:�ߑ������V.��1zߋX)�C�����n4c�PN�T8^�!���1�5�*e�{�J7��nK<��ЪJ?�!O�H�p���F�ؾ��� �"���՝�D�=7@��%���E���,^� ��*��^x&yr�C�l�)��;�y�<���f��*�g�%�������==T7wy�i��K�4{NW�$�<�ߛ%,�'�[�[����o%�5;"�e�C���dҜ��@p��A������|�ҕ�3���$j���p�9�>DmW>��Wp�J>!ڥz/�jNH���T�L��)��`�m��;�v��s��^:_�jC��}3��Z2������_E�C�Y�ԁ/y)�A"���<G�?�ir3�o�IPrjr9 �Y)$����A��,N�A+ Y?[L�ԙ+BQ��L,R8B�β�;-�����3�u���uo��`��;k0����ޗ����|�jiQ���x�>	�	�Rb�SLN�_&+��=�Ľ�f!Q#������Y�PŢΚ�1��<脌��R��N��3�?�rOJDy�}��~��(����1G�K:��C�ۗ��_���c_��`z:��@��xZ�gY1g��d��t�.���� �14�$௷G���hK՜C]�f�t.v��Rw�5}` @�>p?]�g������h��x�뷐QuCGu�� ����:�`4& �c�-�k��Ib�q����O� �m$k�W��ې�uE��
�k����U�nw�XI_��=xά��]�\��ɂ�l\��x�c�Xx� �< b��۽T^E�SsG�]�k�{�L{yք����sj8)��Mz?xec�i[x�nњ>V.*ļ�(�*���&�>#̳6��A����Dχ\;��-�6�d� 鶯u2�=7��UՋݴ�����4��`׽�'*�Ay�U�)���e�H�ƌ$�����!���?��ߝ�;ݙ�ROl��[	�x���4_��;� ~:�ʴ��2�	4tZV|C����w���n�LR���W��;+���v�bO"�ACIE�ǘ�X�`���F���/$P������a�n�OnᅎE'U��zZ�v~�J䄮���1���VD�I�>Г����I���b�E�}[9D��k�qû�_�j�߬{�W��#l�_�_��}\�2���
4�0$len3�Sw��~A��d�*��PĔ����3�l��kQ�֫��Kz-�)u�
Z;�'����5U���I�#�ƉD�f�3�Ո��̾Q��?���d��el��f��ED^%���#�ۋ}5�wl ��
��B�UB 126���R;,�p�i��G㘦��R��jb9]٢���2y�ݘQ\�����Z\$��3X��d&j(��3c��ٻUTg�3�����4�����N��X}���b�3Y3*�`����Ԡ�9��
yIH.U�'p���3�^g��o�����
J`�+A��K�޼��C�64����+~+!֋���?��R�"�"q^>S��=_jW�:m�����uSv��q�'KO��|�&�};�Z�0	3u�T�?�ݳ�	>~=�W�~W����J:���f>����㰎?q��ұ��P �o�͸(�tv�}����n�<A�t�����Rk��;��~/�u��r�t<��/U�#<��y2�Zq�v��[f�Oɥ������ޗki2K��ح劲e'��Yb�鵮u��H��)��nG��\L�A*D?�l�e�R��/����4���$����7�/�=���`wlb*����TQ_K��G����r7��V`7���Q���.(�z���I e?}T�!�����U;5>�����X�f�7΍~���[3v����^nu��vxH<Qs-1Y�
�����:y���A	�t|��Bv�'�ާEC�N ��$�!u�2:$Y�W���
2/<$�t�����מ����iil�Tgy��s�D�Q˞����-� Y�����Дʷ<�g�)���L3T��o�r�6K	>	k\U���m��H<�����!J�Òd�W��A�_U!Q�1i�.u����٠���;QA��zk�M����d��Nf
}'w^�i�"5
�����R���1I��}���'BD|���%<���F=.������T�:B
�����̨*MT�Q4���DC���g�|~�XG����9�^��H�g�J�p�����MGޟ1�z�]Y��*�>���|��i!��"��ȵ�/c(:MQU&��e����6��Yr ,�S�	��V�Cw��n哚xg[0	�����<q��4�X��o��M��G�.�W��i�����o֊ض��:��n�_�K�W�k6۬�&Je�f����ƨ�8��]�c�1,�N�z���3��ΗF56�1N��6�M* �jk}d�zWwsP��p����rX�H v&K��.�I�Q��`)/*�qH]X���S9[�j*�^��D.��c�Kr�n�
�xF��#��`P�'{�#4�J�7	ok�����rm�h����9����$���'rP��x�Μ
��t���_9|w�Wϭjw{ص%�q���U��5��DY#�G\�Ł̀5���8c�,~�N����2
�'<+ۏ�Am$��)��O1��wѥ1������:r5=�+��W1Z� [)+a�y5J��.#�7�'��n`n$?��f���aT���.���st%C�G���g�&8����/�� \X%\R�3_OCh:r�c�u��c{����[v4�X���@&t��h�����w�^���`#c;#	��>��O��|*����*�z��:���������������K ,@���fz�����9'|q�3��s1�w�0̠ u��~��ӚL'���v�5�
�����VmSd0�Y�*5|�k���}�F�}��_�뻚X��m�X���ZJ����z�,�}M�U��6b"Y&��;7휦�qj9����>�� �%Έ�3L�����.���{y���yؓ���׎1&Q9*�Z�A���'Y����cYi��}���R�`�QJ��	[{t��eg<�d�z\�R#(�����15�.TV��7S+Έ��mT{�Z>Q�r=]C:=��Y:cG�ś��h�W7E4����K(�t�T]ge\��E���^�D�4[_���a*qc5p+���]�]& ؖV>�f��K��Pzr~iah�a�z��ґ�z�����)��O��y�c�^��AA\�:~�%�X�9�'����?���B"���.�n,k?G����o�5��4Ѥ�y(��e��C.� |�'ʽ�Z�&�`��=�/(���ƞ����ɢ��~�}8��L�]'�o�b�����φ}6�r��&��ϑ�Mv�YЈeN}Se�$d_Xv(
�_gi�w���sO���V�[1z
"��w_�cf'&����+���w��P�e^Qx隴�(F����F�[� �O����!sy$�qx�>��oqg�����u,қIi�j|��f�]8Q�є�#A������و��2���2|�o�1�}�tu�]�K�k��.�E�DA`oA����[-��
�&���� 9�U"�Cx���$WR�en|#."�B�5���;$ko��-�i�s)�s�� �w���_���*6:�"���{��2L4d���i�:�M�GL�)�v��	���6�)��#W..���r~L<�HnS�O9F�V��A���V���A@D�o����8���I"��~ZJ�h��?�m��&����������=�&��3�����7��^]�&2Wv�'p�� �^'T�i��A����-y�h$��P�u �v�6%N|._x7s&��y8��x�0y�6��\��:>p3�\�=�����dV���g:�~+M�\�i��I`��F�f����@����B
�(��r���s9���'ُ�R�M.�C��j}��j8�n��Z+��������!\NɅ(�k��tVT�63-]�K�~�,�\�Ɲ$�0��#T���V/��n�ن���F40�-=�K�{lD�A�Via���k��h��n�c/�+ZQ���	��'|�.!��t��A��l=��f87�oN�ɪ���R�3�G#�oZ7���m����$�b�>&�����kj�tw��S �#�0y�	(r�*f�Sy�I��h�p�)�53��|'[���{�UF�q�˘�����|��Z�#\�[�<��D����S+���P�>��bt�\�����V�`@Q��gQ�c���C��#�0�_�9���yG
�(yAi��� �{�����ei��duB�V��A%T�B<>�h[c��j��=�w��DR�8���:/'N��ۢƘ�}�h�I���/�*��p�Q�*���z@��ܠiG�	鏣{9�L�����Y�*&�g�u�
sY��ꦐ��YmN�	�΄ۣ�dRD�����lعYfg��f}����'X�:S�>����((�R�t�n�v��k���ݮ�0}"�t����u#<#�h;/�����?�����&]��[|r����r>��B�l��7hM�{ou��u�ʯ
�i�,zG���G��(��z"�.�XD<�R���=}K5 �ӯ�FP�0�
j?UTQ<�m��-F����B���b�vu`��PX�_�hsap�O�i��f��0����s�¨�D(�"�R�UG�U�<C��d�%�f�`>oe����_Z�+ �*g<<��j�l�SXԺ��0�����E�����z�,}C�\2g� �U]�Vd�>˞��J�ѡ�=��/X���,�pb�gG�E'�Q!����� �r'�J��ݖ����*%�.eo��Lv:k���Y��hB\$-��/w�-Pg։����0�t-��� ���� R��ꐦ�h�$	�ãdX�W�L=�=����~(cM�i�{��e���)��֡��"�k	E���e�Y��3.��e�0��Mm���+{��=s��S�񎙀j'�A���wt�w�_��#kt{b�-�'Ȇ5�C��5��팹�~�j��7�~%!�3�d���i�[�Ԕ&�M:�x�@�rP퍙A���3�1�<>�5g$�p9{�ŝeM��U�
��,NKB'4�^���,#���屯��5�aT��w�HL^��Z�u	�7;*YwP@(G�����nl� �i�HmP���C�P���:?��ѳ��#|�I���l�0���*�t��E�<�X*m�i�X3�aK��q�,��0����.Ş��|!5��A��Գ�4�ԌG����m�S�$V�}r%Wr����nO �g��a����2z0�_?�P�Zx^[SH�Dp���E0t��`@�TK�Xt�]��ޞI��e�b�	~?E���@�H�T~_u	85p���>
C��'@GK��9>})
��򸞺֤�Y���CM`'O"fz�����/�����r�(b����Er^�3}p9�n81�uQ�N��Ò(�7��(�	WF�ڀ��y��2�O��r�(��z#i
?Ѫ������s����a�L��3�׮�Xi�"֋;fnCb�Ҧaǽ��E̩a�0�1�Y3�be��B��E�]D��?���X򽊫2+��������4�Y4����s�z���X����	��<L�+�ſ���$�%C�i��u�t�Q�Z�у�Ж�g�8�3�7�8��g��xG�2���z��{������E�<Ü��Ǥ���A�K��'��7��`�<7=��7q��T.O�t[S\�up�աN�Ȓ6���7kic���3�E������.���A!�����)��ĺd���mb��{7i+�D$T�'���k	�h�>Y�ѹ(������IH˰	u�l�/�DN�c���9~���߃ZǞ˴q�<�Ei���[k��h9H�C+��`N%�	Ef��ԱQ�ydZ����i(��Jx�[��C,�^�B��W3�E�#⍹ETF��E�j��z����ξJ��"�Ӫ�� �QPxn?�S�v�e�BN�dM���=>���,����Oz��:���A��|�sD��Y;��[��g�D�&m2�ֳv>7����.��>~������{�n���H\A�5�P��Q~���%�i���+P�e�E��_	�kN1�G���窳}�9�h�Դý�����b��m�����'L�R�(f7�]��o�Q�`�8V^f&2B�R�C�9�0v��Y�^��ξ�h~�P�W29��������=NOp�"��sM�}oQdr �>öv��H�9��6�o�gB�7�Y���l��}e��ƿ�����Km�o5dõ�{���G�������(b��&;�
y�.�u-�#�0�|�	"Êʥ��Kf���+�[����>���wa�>j�-p��K�����SFQ1	J��)�Ő���i��t��ָ�X�u�U�*v�W˹i��h_�����fv ���>3J̹.���M�R��d-�EvZ��a���j��q��H����Îs�u��H����.� ��3�ʱ|�)}L��M6`:J��LZ%0 ���Fҵ�SBF�<��Z5Ly��S�ܵ�T���d�陯mH���v�);k�y���^0�u@x3~�=����d������^c�����l�����@�����5M躝��@�ވ���؉U���YU�Y�V;�e���n�mH�Uq0�|;�#�f�����W28���w�i+ ������t��H���;˂Ts,��W-יL��ۧ�ur�i7�L�_J޶�x���+�9���-�'��t������/U�j᰷�� �[�_㙝αg�3�d;�#w%��������{�
������q����,iE�w�X���V�?�Z��;�� )ڽk���aRx�eᅮ��0���9��"wp//����^2��V2����?���� ;|��*�F �5����u��IFuA��`z�M_�J5j��*ꍋyn�����ߥk�aH�xJ|{����cIk\���fQ
	��+�U���(�*k�[k��1�I{M����a�XA��w�6g:G'r�i�&�`�[짥{ǹ��������<�X+(��Ԃ��1��G�E\�v�}MO�윟�������L1�<b;�q���`��N���j~��:�[Ց8��׵�$ʎ��j�47[8 /�vi�Ͱ����Q6��j�v)�S!�6�����2m�)M2z|-��*J���i!��xz�>�eq�	���`b�R��NR���K;qG���:�	�l�\���V���Y˱-��G�T�}����gE��Ι싓�*�� (��;i�w\u�!J��ܺ���}Y.\���W$���D�r:����+�{����zh��_J�߻Z�*G灟��Y��>�	chG&�Ub�.r�ʌ�Q�]:��o̎�Ϡ�>�z��5�,�Ù��Q��}� S��q�j��Zemc=�k�A���0j���D�k#e1dǅ��b��YP�d�Eإ̺F�Eyd�#l0j�y���\ޗvС��n*YB��rY`��w�w�A�u*-&ޟ��Nˁ͇�T��֌u�jI�B�8v��⋬6X�[�]~��j�Ϣ�N�	���Li����G3k&��N8穱�'����2����.K�h�iR�a���:Z��dזC���q���Ƹs�~��4S��L�U�<�2)u��m��D�77M
�66�^��\X���_�]N'l���o�7a:��uQY��uƁPa�n��h̀�"Z��ʠb1�t����(-������G#�>�{l�\*w,��'6����ՠq����B��º��Q�[{^L6a�ĕ��t���	c����d� �g�qo�If9�U�s÷B����3f3YRk6��!(U��_��R���e�z��}dcF�0���i�陓ZX�C��A�5��nL{p�h0��^,P~�IՂ�f��%��hU~�V��Z޵k�i `�'g�3�縵�{����	#j>�1V#�����(��=�?��N��g�ɉ�B !2�g�M���'�ߊ��Ob\�9δ*�9Pj5,��\�y�	����Q�`���]g���NFin>� ��$m�/anf�2S���F5FN!��L[����W=�� ���+=]�K�6�M���x�Ud�T ���,+h�{S�,���	���i��~7!�Ә�I%���1�Pk�E~Ѽ
L�l�	�J�02�c�)�6�cH��nM�Ċ�[,�O��7li���-A�"�;mbf{@#��,(�g��)���L6ٖ@��	���ɿ��qR� ڷv1�g��+�-'�K��œ����Xs{�_����_ ��A��UsW4F(�`�r#����"��c�@=���Ki�
(��Ix)���UlS�':��4�k4{���?�Ԫ�v�#Uu�O�-���F��A��R[_��ݞr��`a5t���>��6=��A�m (a�����?~�)zô�=8����u�4���O70�@R-��&LWJኜƻ���,H�n=U?�-cC�:�p"���a'g~d���FN�u��on�OV@�DF�R���7MvD���܊p�����j:�3�b]����~-�iz<E��*�\�7��Ҽo�6��+��!
�1����$��I�����2�1��#c���䐡._�.FgPk�ؗ41�Q�{9�QFk����>K�f�Ґ�F������$�^:5�>��L©���a�A���kz1=��sM�~�����.�{ 7�+HMm�����m����?���v��JSAq��B=��-'�1B�����k���9���<���Dpq���!�O��A�@J��c����w�}})�Z��=ឮ|�a˲�z�R�l���mB���d�ݛ*�E/Z7��e��y�zS?�� �C�f
����&C����uU�w?��������o��þd���m/K3�St�m��Ծ�`���>0]��;��C}�dz�t�'�1Zn����A�^�S�Ԏ�K�|)�?�:�����4���}�K��=�K��eY�VKE��̭����w�x}�4IXܤ��Q�M�8�� �N3�ɽj���=:7�X��	���E���3��T��^F�L��c{� #Ġ�8�m�ݰ4��cֈ�-&:�x˟�F��x����a_��_����Ż�~�{}G�&Eԛ;��(AX�T��7�����$��z];S�m�d�7��tI��g��v���2B���pC��s
�;�J�[:a� �;�9���2TNZ�~�us�H�ۛbe���X����XPQ��V �!�i~��3OK��G������C��[@�<�?5�1�;��%;z�2�>�L�᤟��诘�u�Kj��JL�w���h�h"�Q,�W��jZ�:�g�6:t��F�Ϡ�|�-�P΄gn���(6`���<�fx�H,>G�У�S�Wv��� ���!I��o�n�Ҏ����YSA����ڤU0��n	cVY$xW�������Rc��\��%��Y����8�����>�eس?���}�B[�R�x&R�3��ݐ&�M��Er������|�C3��emc����D#YSl�_U�g��#��2����l�(:�@�UNI�A:�>�d�����z�5|���RG��!�	�	cG��4R�[����"E卸}� �"���d'I
b�+!B��M�U��2i���i����#tCp�YɖuH�r}xb�0 �� F.p. �4��ۢ�隚��%�ؕ$ڤX�?��g,:�.q��	b��~*R;c�Z٠ۖ#�($�l�!kb"c�N���إT ɿ��kZW7��oh +[�Qa_��ƀa�/����^�D��{"b+�^R�l��;��m����^i�y�pk���N���H���!�=�a[n�g�^o�@�Y ��S�]�ѫq;8�I��*g4�������u��@��a�2#�~cN��ñ� ���O\��@��5d�4EUQ�aѾ{���yAx��"�Ů���47�4��Sf������^���v�暙S�Y ��*�0�'��t�f��I���({ųV�L��d��p�����RA��}�<�2�~�s�=� 6ɵ���]�>u�
����=]�ǭ�5R�s���w�D�7W+j#�	�K{`g�❱��VhI�1�|E{	�xE�aw��}��-ț'����U!��#8��� ��xX��z#HDw	5zFzpI�"�O�̡{C��"9�-A�>w�`�t07G��듓� ���A����}ʑ`PC;�?{�, 	Q��EnU�RL�XL��"�)�>^y2J�<�~��t�|=���������������R������}�AqK��K�?ky.jg5���\5����L�r��x���G�F�м���o��PA���X֐���~"�׉�/o���-�"r���F��� ���(pln��@�?���R=k��|�|d�b?_q>��{�m�ƺ���]#S�i <�X򗟟ؓ��c�y������5�� �������luOp�-a�	�XE�4���,X�
Ko�POJf�p�A��69���#���#���Aֿ���������y�?���*%i�����y��=g!��[�\�A��Hxj��m.�_��-W|�����d{9vZ��?��ٕ?DU$� g?߶2
��꽮P���|2L��*w�O�:�if�h�.i]��1�uI���l�aNz�uהra�S��jr<�:�sL��&��X���0�w�_��7dЊ ��yEV�$6�]�+�����s�˩��:i��G���=G���*�"y��6l�/wgg��<���zN��lNɶ0H���V'A�zP�b���R�2�R���3�_F��5/G�;�b�.���[:��u/(��E� �<�_��1۬E���N����T͵��
<���j�o��*⾄4��ip[�+Y �i
f�,b3w0��:�a*;���F�̈́Ud�
�Lb�����N|�1�`�*��ИMJ�ք��r��/�c��]vM|�&)6Ԁ�j�r��ʮ@�e��*v����~��!H|62��U�Hp���(���D{+.'�1c,���q0B������SU���$��Xʢ͖����	`�SP(=i�^5�m�:���W
�)���j�4}��.�C��w����t"�K̓`�ȷ<Ŀ�PȨ)[��P]���;�P}�+^��Z#�}��<,)gZ�w�-��JL�-[i?ZqG����P�P>�b�v�u<����6kd�ԑ��?|����gNl��u ��^a��IS��1�3�])m�m\QwCRC�5��eS�k�.���\J��>��u?�	ť�C��E��COo��]��^��b36rP��`[YcJh\���!ux	�F cV�����
h���#�ڇ�kx@��p���;|����5o���;�/U6���bH���ow�{a��6r&E���n�y]?9����a>w�ɍ�(S��w��O3Z��} ����On����L��t��V:���h`��J�n ��?Ұ�ҀQLX�R�i<�wk��M�"�#vTad'�0��s�H�ZE�f-���'M�B폦F��uݎ�'V�.+q�����吧�s�(�f�<�(�9���@�����Vx&5��լ�|���.�h���x`W~����Œf;�	��T�Q̏�"�GL
�m; �|�A�Y���ӑ����$����R�a��'�/�昗����O��@���a�ɢ8�:��dቢ��E�+�U����x���,�.$D���c`B�|ԝP���a94`}�\�/��ǭ�|�@��.Q>��&�Fa0�j����+r˔�B`�K�F|��<t�89۷n�S�D1Ե��(��Q��L�Q1T��2x�޳ ��W2y�V9(��-#8�oV��c\JM�K�v-�>�9B�W�0� ��b0�z�E��G��3ȹ�3��.u����"
0��>8��k_x���0�r*�@X��p����>�a�� 	4����)���
�cU�m(J�W��1R$o�[Df�./�4�$t�|���:%�Zs���$��	Xz۰�����v����3Iri`��(F0m���{�˜�30�=NM�4%�����D�\k8|���TM�";AdUuO�Zƿ"�<V���`��Ĕ�P�x8޳Sk�qj��Oˀ��|�t��j�����;�X�yr+# yA��y5�����vK�h�.��34�rQn�}�lg�}���_���H<���Kg�O.��Q���ӔDr�2�IfGN���~�z�E�l�Y�9�k��ȶ>�5(P]!��9)�b]c�.�)��d�S�T�(���SڗDgV�ir ���Fm��aBvC�u���a�|�
lv�:l��19� )G��̝֔r����c'f'u^zG��Q�Re�~Y���f��iWo	e� �*��~�p=o���[Ȟ!.K���.�'${0pAl�H$P�&���M��:]׿�%&% ����8���k�a�H��9^4�V�j��&X+��7Y|��q�D���_"мQ����ن��#Hs�Ё+銞���b�AH/����c���s��2�~�C�����:��
����]c�H.��Zj0��G��.o���|x�e���v�m�	*�	ŰLոm�1T�Ż�⽶_���:!,�[���:��� -��c'V�)'���^�-9����ʱ���Dy��/���٦#��X���Iy�:��='D$b�>�*0�cy�U~�
��m̒w	�s�0�z^Y��c����a�_��R|L�m����=�z�_�X��]
ܮz��m���p!���m�!�@~Y�������1�8S�D?S2��1��ċ�0eF�Gu4��qB�J�e���[��VS#
���P"ۦ�j���Vi"���z	��jiW���!�W�/��b��"����fJ{" �F�	nYZւ��v�D�pfNN�J6D~����NlN2)'��L���F���3=X/��TI��3�ۮ������m%FܧZ���2�!��M#;���s5�/��v9�[�ϱV/���k�/d���H߹f��Vfnd+�%������������h���+�pr��i{>/;/�`��59�d�]��d���UZ��J8
� M�@^��J��7�"n��/���Mɋg��s�C�b&�����5����~0R�L�U^!�j��x�Ц	W���b�J�¡�^x�ll�"�z�r��(2d�ذ�:��g��ۯQ\�;��L���Y��?x9�&9!�,9۟D�B죿Yy�޾>"��&*�)}�09Tmv�ԓ��<�׿��|�\�o�jK1�_I�Z1@ڧ��D��;y0���>|�4#`dխ�Am�\�1y
���/�:�/��*�v����`>�i����.3[)B1���9p����0N�lV�$��'R��~LQ��z�gs��_��ء+rM�2�2�����a��8�$�0(j�����ç�����b�z%m�!�D�^�G�5�'J�jj� (<�9��=�����Y6ҹ��dj��-�O)o�)�ì��XC����-~�ܔ����LT��T�E�����yf+̚����ٕ��f��8<nJ\�S��"Їj���96�������sgIKrf�aq}�D�ς���E���/�_V���  X	%��(�^�u���1l����Pp�T����zUK��2���dKa�`�}9i%�P�37ӫ(Q!5*��ñX���
\iC��"�-��"�8X�dҲd{�n ����(��g�o~������:i��^q�W�S��� ��w��n��j�bk�NBx���@8�]��S��%�5�E�O�o�G��*$�}�������l��>2�	-��Z#jD��W�3��!PU
&[������b���a�pf��Z��Kx�+�؍�u�C��K%�:$��cs�������О�qZ\��POO1�,�*`C����p#v���a��>_f�� 5*�z����h8c��E��Y|�&�Ɋ�,�?%M��Tgma��x������h��	�s�!kp����ͽ�n0��`�7���k��,���N
b���ֿЙg���!a�f��}B�E����@(�8��_�UPϤ�{s��^�P��� ]���.�9%�n{_pέ0�CPc�	��� ��� �f^#���_Fm�s9Z��B�3�P\�� Z��gр�<	9O�B�_��p�4`�f���h�Ɉk�Zt�WRRJ�q�s���B8�	�8�`A�S2a"��1�R,x�+��)H�>��ga��[S߇Tw|�i����Sa�l��JkFH��}e��lof&셵�{�Q��X�ZP��7�Y�)��nA)��6��	n�T�#鳼���?,P��!�sZ��������s3?S2����MVf�UO����īCo�B� ��le/em;1K��G��הϿ@���Қ����XM��ry`��t��7���;m��g#-��D_�U��_�}�L�����>�-������H�3���s(�0��a��=�]���u�Z}�Km�֭��ʻU�xi���d�qC%�3&y�I���-k�@�b��k�7�W�C�~�� Ll�%M�y@���x�V�h�iĪᨰ��BwvZ�[I,*4�N�_�cr)��M��
�/�����;5��ƶs�7�mn�"ht_͵4��>�4�l��~EXW2^��z�'�ݠ1Q~�׿}��G�Z>x��Ԇ�^H�b�g��QD���섁�O��e��+�f�O��r��y\J���Y(�����(2��d���;	KaCD����
�� 8���\u��96��3iC�H��3�jR�Aۉe���M��@�����h�+���tr�^SQ���:���X���6E�7��9�����j�O���[$�1$x�5�oj�����f��>�W^�M M�(��m��a<�����,���-4��|��9�S@{
J;�8CV�j2�����0VH��A�&H��A���ϛ����\�A�#y��c�d�X(��5Qݧ$�q�,+�>�Z�o_�U]+1�n�����e�;�~�0�'/���2���m��v��ùRg�*�����Y���i�jVyi��(,��X<�ԟ��R�|��%f�'Q��y�]�O"�ܯr���'�9�⤮�Ȁ�Ls��0�d,M[��;�j�������rK�8���ۥ�	Nj� �y���I�W��+G�Q�}�Iȇ�g�jjC��J��&I��A�����E}�L�$�d�NوP=0s�8��-��D��v�o�D�ևr�����'��~���'�8��W�,Eg���$6�<~hz����Bv��F)�ـ���87�(q�����X�
ݭZ��A�ΣY繅��!1x�<���#D��
y��ώ.@�IT�)Ű�ҸP�3�^�j%�������4T�����^�m����o�F�)\ �*D�o�2�c'����Q�u�� ��]pa�<	Ir�s����Ka�������cX4{�OR�>��Զ��^"gW��u�WsK���o`�Sڞ��#֤6��� h�8 q��|�4�/�4
m�)�J$���Ä�g�����e�tu<���,�C��F�>dm�[�����i?���@6�h���zg��D�Q����5���G	�xu���S7
�q���dp寜�6lLB����Xݺ�ߍ�W��1<��M�Y��>V1�خ�nN�3���Y�]���%=�*Ni���hk�4� E�2xa"�EI��3���5C�Π�/����H��#�fU��u���R���l����#��$��t����U��8�N��Z77���_����Q�p| ã7������k�e@ɓ�-ۄU�����CV���4�0p{*zEU�|�����p��O�q�����XN)g�~9[�7�l�^~�
�3�,�覌,���
�*�F��r�y��ޏ��8
�H�G|�����^ AW@qQ(ޭJ����;�������߇�t.4�o�̘��M�3l�M�#t����a�U�/b�!��~\]�5M��>�n����9`���I#��7��N��5�AQfi	ǔo0Sj��eܶ������_�yp佊@!%!	�"��@! �2�� �w�GE�_����$½W���5�3uF���nC|�O���Fe��T^��O. *�iC�ej����qL�?ǜ���6��={ċI�������BX����+�e�����R D�,o����+S����4��c��s�̇( ��,��'��$Z���T܇�����<{�Z�cdQK��JT�#P����"E*�N�]*��@ep��@>��1cu9'�a���])�m{r�jD}2,�n���;ƵB��z�A�4��y�ii�G>EL��Y���9cĮ��*v��Y�@��6PFq�	[����zF1O��������>Y�I��oF$ӽ�z;Vy�g�D����.�Q})'�-�$�f������HwcW���0}��^�x�-�Y��0P��"�V�
��x��SQ4u0�s�۬�Y��O�y����b_�l��׉�<�('#ɳ>8�\&y",z�u�e�l`��'�9A���Y�j] ��X�N����IF'��2�V�.i籲�Xn�k�A6�GչrW��X�!�3���&i�����D�����]7��Ny�n%]H;��@�T���zg���E^�6h~��Qb�8��t�~�ϓ�qj+�?�����L��H��#����CPb��=Eh��n���ŵ���"5���_QI�G�G��vI�p'�s*z<;���I'G���Z�l`���b߻�C�mV���jp0 �r�%ng2v���o���j�ˁ�[��5DH<V��~%p�ͷP��: �K��ۊG7<�}�����)_`��3OG�� ٛN�V�l>7eȄ',Qjh�1A�Ĳ�I˰^�D�e6ۣ���}l��G�
��g�e�?���%^oT�LWc@ɘ|�uZp#py��E��֚�62�~�ZvzxK3�:� ǪO���<���u��iѻ���G,k�����`�M���"��d��
�O��͆�P�4����	>ei{ԺQ�iI�S��k��:��d�\AU�2OK&\/I��r����]YY�T,.n�lE������@�v����`�=a�	��� Y-�M���3�Z6 �E��c���[>G�?�l�ډ�sp<k\��@5�uƤ7�L�5�;C`�[۱`[G3����x��؜�>L�������K����w���N����\q�Zz�<�-��?��ș��,� ��`�r�(��s��z��q�m�c�h����\w�N˒k@�p�1q�cE5���l͠�\ی���<�K
 z�A�֙��N/���Sܼ�6�]�)�@�UIU��lO�pC�?w���{����;|x���xt��C5z?U�a��`=��%E��!��	SN��
�h���/,��ԶtG�h�]���+P��{D��5ɴ����
�O7�~�+������_�kEK>�N@s����o�
*�6�jZ���f�^ϱ+�+R�E��n�`�W��|�hG�,wuB�X?B���UH>�cX��7�(�������k(UE���X��m^oRj�%�_9L�b��쓓-C;kYЫ���v%����P�op��>�T�%��)�X�����|.陵���@�-�DŏB��`�����.�b�-��Q�;8�B�������"L��l�{Q�{*�4��hQ�Z؅O��U��MDP^_��|K?�!煆ϋ!�L|� :�B�	��h|5�@bb$icR&��rpO�K�V���X/
�y�+.��̟��Ӓ�P�]�����[�$?�s=陂�M�De��Q�ݷ=�����6HFCm�7���_��<��LE>�:�z	���6B��"��$�����Q��y=������-a98ڕsF�ĺ��5��u��LO��(��.FpP���Q(2S��2B�+%��G��=�:6�c��amLYP�0b�º�'h��
��C@�d�������ب�G�V��#s3�1��l4n��>�u N����F���{���;}�G!�M�8qaչ��A�/�f`a�ȣF�����)A�Ǒ[f�>�SD���Z$����ԋq	�(���2"&���(ιM�����B;���Ƶ�Y:
��T�ܸ��=%�|���(���t/]z����ժb���SO��k�zgF�sS.뗨�����?ݘ�r��;8\u�����mxy�iv8_���ji��&(�ó��D)�ϴ�BAG����6������o�'@��1(2}�� ��ɬ#��$�������Kq�%�]G�'t͉�*�or�;Y��bW�ĉ�,�	 +�F:�`!i7Q�8��?�[��#.Y�Ϙ�������6/��9
n��(�pAn����䫸H�gS9tLh&�
�x�����5�#���2�'�+���OP���G��p?��߻h�j���F3���D��|~�ڬ"��ײ�sÇѽ�^@�C�C�~��Ƅj��}%Cߊ�����h�_<'���k�(�0�?�g�Vs��Y������[��?�yC�Y���|캆W�V*����կ�"6����~ �����TQ�
�\���"�s6U�yWHF�ԁ�(�J����ؒ.��g�.�%zv���+*Z���{q��� ���+%�W��35'X��s�NZ��%qBA�;8'sg^o8A�6Ѷ�ү��:Z5�i��
l�B1i�# ���^R_s�<�>�)�4^���Ĵ��UAO/�3|h=i�N2�d�g�#�����\�?��ҽ���[}�.z�3�Ktc<P��+����9���س��
$; ��e�c�+Ø`J/�?_P䫵;�
j�R��>:ϕYd���&f��*̪�;Gr�#�{�f��&�W�&=2i�8� 4�#=���fϋ��8�!��e�}������E�N��Mtܫ%���5$<������c7�`�[k�c�]��/�{:^�{���6/������Z�3v�>���!Z�r%�2��[�jϳ�ި�(C1!�l�/��y	�J F�j���N;u�
��i!F��	�)p�������~∰�`jGKA:X�D]۫N�Ǖ3�-�3ϸ��ݒ�e�
]Q�
���$z�
tH�NgTA�r�4񳮃�:�3��g0�7�_9=Ï������.#E�����C��XD��W�y���j�kf��̕Κ?!��iB(U?k@�'����f	���ɞ7���(d����Sf'��������C0� 9&�C�������3��*ҵA�=$�D��pt)L���g8�]��Lg |M(au���D����/��Q�(�K,��(*��ﱂW�����"a�$��[��xw��d�:i3��ÿI��0B���?�G�߈\T'�c���U�.4��܂����ށj�Ҧі���%k�~Z�u���5a��:�4���P�-m�΂� ����=>�$���%��惱<
ķ�'߼i`�F0ƧZ�#�ذ ��{���\��n��^��{O]��K��]q��]fXK�i�>x��~=�T�d���n;ߖr�E�,եq�u�eɞ�.����:����6��Gy���a+�HO��4�P�"g�c�y�d>R��<�\�	���L�m��*�����������Bk���ѬE�OQC���WO�����DZ�2��#�췭����Ʈ4Z=FO�����4��Rw�7=�_��������I3���v���ڲeL�א0���c��wH��J����no29���G�+����p�O�&�Cl��w �|��`Pqw�RSj>:I�����
̼� �yb�D�ō;G�<�dBR���M�R�
gI�Z"�m_y��?�063��w*m�2>G�{D�$�c��^�Nj1�ε�b��2����H�;4~���0��";u�sa��G�G~a���~E�?d�g�y5��S�a]&=t����.��z5B�F�`����@s*ۖ��S����_R�4��/�Y�#�]��4�l�pW������e(�깤ׁ�����iB��9��SwM��?�8��m�sgɹ|��p.�rU*����Ù���q��ZJ�p}���ә؍iV��ɭԳs?0��Tov5sD:���r__�{�h5��)R&��E�n�!9�J�]�fC6!��"�.���ș��p�.��U��p��W�'�B�Ҡ]l?2��8a��vW�~�O����C���]�61 �v�4:��;��ϥK�n-b�Lj�+��3N{�q^���c��ɬ���x��&�_7�U�AVq���pȴ?�k�o���Z�skf�F+ T����e�N3��YH���xۜzε������Ԣ�n���}�� �N�����*c���-�$>�AŰ�E��1+��W[kv��=>xs�?�E�!�9s�9���0���޸5W�8��4r^�
U�i�E�X^��a
b#?>R���>�zؿ����f4Es����]a{nxO[b�.���t�%ØZ���'d� ����;qNV�N�y鷪�~<>�`s��;��N�R��N�YK"dG֟�#��o�^�)Z�B��b�l��6�?A�׍.8�����?��}e�sΝ^e��5��{��mF7�"ǣ�Y���"���!*|�䳘��|�Y���L8�F:�oaX�G8ک�
D�����9&�}Q�權ڄbmh�?p�F �����͛��`��M%Y-�˳�P������P��T{Q� ~��2�b�H(J�Q�^��Q�\'��$:���>�+K����l;��#u��F�ǯ�)Ľ��s�B��ؼ��VT�A���t���t���n��;�t�kH���;A_�NDe�d!�Z�7�Ro���!0�1��źX�'�ڨ���#':�"�s�,�;�P�-?�],�z�N��ǁ���a�Q��2�G�I��p���<3��-�l�ӌ��ZUR~�v����O��u,PE�6�3�i�y� :"clP8.�� ��6�Le�7�g���d1�t�m�8��*�)�W��6n�$x���O�,�	��|�6j��斥C B�����]���b�C�܍Ⱦ�������-���{�N�j\']=)�B��Y�j|�qcQܛ������E�ՌD�ib��f�Ϻ1)���42a�_�>���0CN�-�mcEx0ѐ�@��X^艟s��xH�iG�(�,�SG�ِhd�M)*ٳ�����^���� �����w�V\�tp���2LC���r�D�qIc�:��ɻ�����͈�i��^�#0!�	��Xh?f=$$g[k�n_�W�J��n��wuɟPjO��KΓ���v8���j�!��QW3Ǉ�����?�V����`g!�+�q�Ҡ�r�����楯_�?pn�RL���Mq�ׇ��D��捉�8(V���ct��"r�����4Y�L���{G�@V�`��/��0�U���h�(�/�a���yHy�7�Un{MFGfO�Q2�򁒧��u��!42÷3��1O/�)}����@����XՄz�F��3a#������T�תyt�F4,�
� ��J�`��r�mJA}O/��M���b��ȱ�C�W�.�ʛ�'��5���b}��
T}���H�+��\K��F>;�_v��ekݹX�uƊy��=+.:�7b7B�A�e�$|4���bq<�٢Q��5��Z�߹\\�	�C���C��:3���j����(�7F3�P�/�����K~��~Ldy3��u�ow[����e"d��yY�i�I�YN��A��:x]�щ*�e8���U0�������
BX �D[ȭ8��3�<"��{��
�$ ��!�9,�����n�����ML�0d���v�~##~�������"�TC�;W����O�����4��i������q�����j:��3�>S��b��62�NV�ش�r�;+0T8d�Aw2��Z"�k�RV� �����d?S�?�y�9l)��V��Q�t�-u載G����r0��F����}����{�U���-K�F�i��	(�d+ړ!��t{��'b&)i2,�o���qj�!����T�NR ��_����N`ݡm�9��u1����짦��QW��K���[�����{�,͟t��d��@����'K]�U�|�YNF<�`��<Ef�pթcN�{E�K��1�2 27]iaO��t�>cx��9S`���l�:�tӂ�ԍ1����gr3]��n���d�o�#H"��������'5��S��q�`�-Ղ)�LX]	���	3y�>ʹj�_�n0�U/B7VFWƃ���?(�;	��+}��I/؛<�6z��3���=
���H�n�����K&ms��y\��>fC���O,e��>԰�?
;ʳ��,;���"��Z>E*�Lѿ�tHr	l�{�jh���zy�6C�堬�bH���e8Q#ai���6gR�D��c�!rf���@��������kax|�OB��2z}����6�z���[�:T�z��ˉ�6%�&%�=�]&�'Pj��ڒ�;W��a�ױQxB��L����&���98 z�Qs̠a��oǨ��"��.���4)]8_�����V�	�0�Tg�S���5# .�6Ή��u��;y��r_�(�nM�ݏ�2�`v��|�TU���~�)18����qs��o����Aſ��3��)!��^B�o�ƀo#uY�aF'�8��8n!^�$�9�Rx�8�L�3�}��ѮRg��ɬՙL�t3A�һ�"��-N�wK�;��-��i���纶Hk`�d�T�]fS[ŉ֨ĸ�����b�����w�'�(��ÿ��W�ׅ�ZUU�4�e)������+H�T����8���4����&�X,9sc��X��2L/�'��)�5G�2Aw���U"��i�-R����n�K^����Hl���]O�UKU-�8�_�H}�1���q1�]XS5�T�Y@��n�P7�`�e�Bk��� �ʒ����Q�g�@��9�,�{��Hi�-�dy���D�8E�DG
拥c�ު끋�lz����&��=���v\�~������r��hi�9����n���w�h�-)vߟ�!����+�T��[9U&� �9]��%1�Nm��m�U�a*k�ZM��*A�2����.kD��?���|8i.�p�;$�#�����Y��m�m�A�H'����oL��8� ��yX�3�u<�X�N_����=�#rj���}uY�(�Qї���VI/:��4��0�M8j�3������B@��4��^�b��a��`�P�)[5�n�w�I%��k�R�qU/P��ؿ��M�G$R�P��e�W�+B�����Ƚz�T���F�U�h��5ݼSs�d��k&N�1�,�=ܯ����,��cE���͏#�~ħ�����
LaL��O�9�-�uK'Ѫ�#�C��4'� ���˖B(��L�7/���g ���NL�-L�dE�1��d�/s����`��z��`�e3�*d�u�T�A�*�#��#�me�ń�;���t����������(ͳV�[dWɂ�x�G�%ˋj��$�T��k�U���PH�;��K����/�X�Yg��E��ȶ���Y������@���d���V���F��G�^JX��P�ٲ-����_�#Dԍ�\�o�zji�P<��FZ�sC���=��8т�qwAbџ�뻤�u���%i���c�wRs�$n��0W�t���g%%�f	q�����[�pI[���ݼ�R�>	Q�+�#f7����U<�����񻪀�Ǔl��3hE��W'?2ڎ�cjj��S��x�2�[tθ%�:^P��o������/�wQ!w�G���d�.o��
��T�q�t�e�N��^Z/�'�ڄ���E����qR����=��$eS̜�Ln>V�p�N��\(+��5k���j�ԉ�������Gcn�6�D_�I��6~�Y]3�����a��8.�MIJ���D�r�/ޑAP��{֋����bz~�ψ��� I��A�8���b��OA7�i�*b�䳥����2T$�x��r~���coUt�3��z��L~|�������~��qW��e��ǻ���I����d��gr���g�k(�<��\�n皳��O��߇o��Ԛ�Z�s������n��Y�/�R#<[5~�Da͕���ʅ��R:8�%��`K��+yh���ڝG(�'Bi���Q
[ٖ�4������[X���)���T;,R�<������<�N^�K���1��)�r/�+!)��bͿ^|d@0ب#��dJ� EWʰc
[\ӈ��8�R����k��ĈZ�|��3�u��9�0C̓@|�!�x�Z�K)���;�*�Pm[���<������7�g���2٘�I���:3� �)�l��a��Ԧ�̂��^�`��V��-c�>N�4�P�	�[��Yi�b�� PᄜՊ���Q�]G'�L�!e�X&a�)3ק��/�B��x8� Md�p��q����Jc�X^{Y�|���Vs�����U��/s�2�d��+.~�-K�JM+�&�G�|;\r�?e���>0���4{$�������_�̸U��E>fؘ̮��nI�APֵ\
���������0ox���tB�a���)M:�������Y[Fm�j'�˦�._�O���GR���oM���&�#�/d�+��0��z߮�]A��o|�G�Կ��p�+���a9��I�E�@��S��V��@�pd���l���Ӡ�� ��4�&L�����r����1��&�C�16��hs�|�G͸�8SV>d��q7�a��;�{.QY�u�л>��#$�}h��xL3 곋�g!r��|�"�9y�	Ѣw�~�d��3�+�`Gd\��,y����,��(g�ι��������{�RX'r�h�m,�&������h�mkb�vVJYI�g�4�GM�f��U�Ȍ�i�a	X�Kʋ�J��mB�ںnS�14��|~�mA�KvO�6�YEJaQ�fHz��o��q�S��N�b^�t�j��u�.��������x�~�j�3��RX�����O�ж���\��X	�oч�gN��U$ϛ��$��ﱫ*���
9?ˏ����@��](����{���Ԥ;1���Ӊ��sk�Z�V�J��Hg���Ŏ�O�d\���T}ق3!�`�NC����q�+���#k��C�9b��j8�`�j\� ̌P��BG ���鎿����`�<ћ�� ��E���A�p�P���eq��$^wY2��9puMNЍp��{��^)�G�9�����4����L���yiɱ*�)j�amA�Օ~So��������֭��`4�7�15�����N�&��93-B��G���X� }��_BB��c�~����A�g�2�(�v�T)�uQ����욜��Ko�Rrp.H��D��e��B�����C�_��hi�ٲ�ľ.>8��m�mQ�P���vwHA
��\勽����wa�izw�`��8��Ü0��qu�׽�(
{Z��%h�0���d�Vڃ�����%��L ���|u��yR�]�t�6��e�07D�L���҅��@�S�V�]�6�kx����:�vQV��K?J�������2法�Z���2� ��L)�HY�O�l`& �t�}���|�� ��D��^σ��aZ�濢?��	�wN��������������H��eU&��S��&E�<�$�ݽy�ĸ$�As�!���Y�!ysb� B�H�>��!�p�~�{��w������0�d���{�	�+5opn>E�V���y�k�c�	w�ԟƣh\�m������c��>��jK���J�hl�^=���1*<�������� :$P�v���As�8y��b��Y��d��T^�kr��~V�:6�)�|?7#��� ҃a��Ϳs/�@39�fO�l���E�'�`󔁖�a��Zf���n��)z?8��2�R����[�UҮ]����'١B	��	� �Y�v�^�^��C[.O���X��1>C%�/���L�l�ף5TH4A a����?4�hD�_�#���e���1��R ��o���$�zsfFK\�l��Fϻ��h�OaM1�_�~��E����F�=h�;s�.�_�pw�j-�6��Y�/��	'd8�>#󚯠�GH�Ch|��zd=/_]a��%s�S�mk
&_3�3sU��fN�:\���g >c�(��*��+
y�~D�g�q�ط>{�#5e�ZTD��sz}X�x���dpݔ+�/k-�D-!HOH��у$��H<W`R[���)WA�AF8�6�Zt�]㤪#�\��~��6������Aw�#E��=�F��������R���w$����i�`m���N�����k�T	@�Rqp��[<�������t�����r�JBL�Y�I�C�pf��s�FN(f[�F�1�(�h��=@juU}@�����t�����	WN�8��5�-#�Ɔ���������@%��4�/�s�dB1�l-�A(�-��)g9~��r��L�)Hs���p2�^�o-�����ɲ#gz@D.��ޝ���?_;(:����q��Bw(��VsX������[�g��J���9��WI���}F�����'��0Ŝ)g�~�?����%į�~N�R�k� �%kmGŽ0�E�s4ke��ʲTX��RE���ƚ��c�I�@+г�������i�g�՘�Ϡ�zؚ��厨�<�O$0�U��7 ^a��3��1mn��K����*�/T:)�e	�c�c��;(OG"�����TW��բ�����
:�L~�w�B`�/��8g�%f�эunGy%8Qy���i�/�&�wC7 1,���܂De�����$�s���m����vEV���S?�|�vk�Z��X>RՃTfڠ�ؗO�Q3[��V�r~�k ��������t��B��1�}�V�bk�@�1�UƇ��M��5��,�ƫ��Lv˫����J ���
���v��O7��HK1����t�R��i�ʿ:{�\�՛|$z-�?�/�p���͍��W�Cd��5:�d�{M��й�;�/!�]���2� 5:�#�݋ј��Ǥ�����Aae�c��3�OY�wu�h{*B#�gh9, ��b��@�?EE���<�E�̒ĩ�3|���ڣg�:$~�/W����ê>4� �ȕW�JO�%*a��Ki��r���K�a�|�Yk1f1�"����3C�����5�Ά���Zţy���E� D�~a=�8��0�G�¨��:$���D~��a��=g��<�\*���lt��}×�k�� q�����^���^����^��ݡo6#�sEN%��;W�WAS3H��j�V�����qdyl����'�&	P�HR��J+��ȝ�:���#��D�����-X�ioK�6��|q���9Bӿt(��~Ⱥ�Un�yd�H��X���gŨXΧUŴ.��o�1��)seg���I@����g^N��{�2\z�a�&��?G��Y6��k��`��#���#7�yA�Y�����A"<��U��'�!E�:��Y�@EAD�E0,�*e��~��*X@A�D�`w��+�:�Ug,���Gj����#�d^�86�w��Β%�ܿx�=#W{=맬������q���d�4�p�s#VͽD�p�wԸ�c}S���G�q�۳����-�5�\T+ }P+��T�)��M��u�{�PS�|@�7�&��'�vh���4���[�.ͧ�4"���	��i����G�YO����D����S�"$?x�/8t��m�g{:(qz�YǺ0W���
119��ꔷL(M�f�qhq��68��k���&7,8E$"E)JwD��p�˚�v m����B���ҍ2�//d}�����g�ܫ��D��^ٙd,{<���	����=��^;(9��GZ�y�ˎ�h}U�.�L�;�w/�d��j�j���xEY�ͤ�r�h�:H�)��:a�ڒ�����]��GD4=���u�V�[�����}�lN�X���� �P㋎���éP�(>CmU�Ox�p�R&�Y�&�BG�'Bm�0Z���腹����{����,fB/3-n��:ǔ�����r.�}q��')T���|��Ǯ�T*%�,���21�Ӗ��|ai�#�x�;e
�RO��ܖ�-�	QĞ4|��73i�߀爫w��vm��0Z�`	�rY�;�����B!�j�b�[�M���c��m]h���%�n�=X�|�&rM�|q�O;P�_�Y�B�jw[5�]�D�g3LCvr��жe�2M�da�Z�։�M7�N+�pB3����۟�,�h��]���&�t�@�, \�o2ﴞEZԺ �忢J����>��1�O�ߟ`�{���%�<��*QO,�jt�hPz�����v�Ҫ�RF 2�������=7a��5�l��	�ް����c�i���w^�	�2�|��F�,�RA�U���^�2�s�zi���/��]�!�Y� ��cW��1OG�6��.2�N0+Z��Y�z�����Jcd)!�L�<)ۦsbY�W3cYS-8i�9ɧ�Q)�]<*�:���;w�;����2	�z�Ї�@[���H��� ��5�U}`'Y*��"����uʥ�z�P�x�vm?�Hq�O�E��.W�1I`Xh �.P��\$��A=�Uw f�g!5ۍ�0ɮ2i��+@�Wvc�Bهt�_]�M�hEabp�+H̔x���lc �G���$�T���z� ��	2��tv��W�Zv*�����o>���8lɏQ��{F��_8�D��)��hNۥTpi���N��x�S%`�'�7Hjc?�+b�=�E,p���M>]؅�d���	:�?2����k�}:�x����#kj�%�m?`@*���PRi3R�qk$��?�w���ҡ2���5M{�9�\:��s��r���/=]	>���$Nq����S��7sIR5/�}<}{��,�U�xd�L�G��|�o",MPut�di�uO���;J������*2��}��/����x������~/Q|֎=�%�������Hui���QQ����u�ҕƽ��&�9U�Hr��R�w�kU^�`sb�%�@�b�{���Ԃ,�S���,T���ު�p�h���q9��1Sފ`[��K��Q8%~գ�;�Y�T�@iv�
�\K���t���Ebڔ�j�M^�lI@��<�d�
���uy�8�'$���/y{3xA� z$LK�Oi�$�kB��m�8��r�ڶO��c��R�;tx?!v&'�Uw�\�����8��Z/�SP�Xd�C��+�gaI�|:74{��Բau�X?�����z,��ϑP��-wc��.�a�'��@�_V�Ns�XA
�Zns�-�R�Ġ9~-�	�:�~�W�p��]pPrkG�i��%?"������$���ߔ/�cg���1���+Z_~B��J5XE���}ü�b��Z`�׭Sd�Le)M�s�&W��,����ng�@��i����7�����*j���WΩV��:��d��:��L��M���v�H�9�����\ZJ��/t{���9UW�`{� �F]�N���C-�N,-�JK@���gU*��+�u�~�Q��}ˡ��\\�&��^7���V<�a�����m�tlϴ#Ws^h���*"ݎ�7>���Ahբ���r	� >P��I5,+d�'ץ�gN��%H��E]�]ty�yh .l��)�L��H�����g_�����Ӱ::��U*���Z��W;A+3� ��&�,�r���0ү|^b��p��8`�9"�f5z�閠O�;�v�D�%V�B�Ge��އp|Q���H���4��s5��x�ЌS����^�9���f/�3&rp^�q����$�ĉ�M��6�f���b� W�GB�>p|U8��ydܯ{��qV���z�Z����!��O8���ɓ����v2�`o5�B��5��z"�����i�����p kR������ۙ��R����$�i&M�u�^3�+��7RrFH�� ��Ѕ�����Je?l�|F�9Kh5nhI��A��.y�h	�'v�Y���b�R���D�
EA�����h#
�.*�A6�v���i.��ԣ�-���  �S�
�`Y�gj��ڐ�!�0��kFw�w0م)5>L^�ά/0�ں+V<˃��23��{��PM#�o4Ѭ4I�	z>�1{M7�*�;�&*�܌��.\b�`t���3 �U��7����
����'�F��>�)�������&L�#Px�p�9pn�l[W�>�.I��O _��$�8�A�1iO7�8IM�f�;��ә�KA���M�]md�.�z�àA�����@�RP��]󙑑H}7y��Gv��!���Y ��9|�"�Џ��/�$9]�M7<��<��;�y5� ���c�]��v�çRc���s#�!p���{%4GM̠AU��m\��I��r�͆�k���6������k*$0������:B��>q7Э��4�!1��/�2��ށ�Cʽ0\v�,Y�x�A��H:��� HRٗC<?<'s8�����l6��ѩ7�N����F-?�d0Yq�DI>&��P) k=E���n�±���3���L���Ə��<��V����`<ذ=��2
,�%�Ӽ�5?ʊ�!"��Ύ
�_cG�����T$I$�s=E�F�Ա~���(�^�us&�p|�"�q���0�J��
��qp�;[qp�a�j轍�@������e	%+Y��l����<�h9F�P�Z�`q{%�� �����ON�/�V�ʐ�?��%o]D7��Wb��͚֒4(7U��H�cg����.���˪ert��[s|v�yz�=�H����7������L��5R��[�i�E�/Z�]���q{04���޲nS��齵"���nl�Q��r@�1��m֒Wr��З<�%�OR9V�QHB4O��	o>ܵ�^p=��[�XvlNm��q��lr�p{k�T(�g9rnCDK�f�Ñ߰��ba=9o�1�����S�'�F���fd��+�.e�&! �:��`��|v`̔��ݪm_��{Ҧ�5i��$T/�M�\����J�)�rS���3���V�EN�F�W�j
I����@A�!9��J#��$��|Y!���(��]�����;����8�ϝ�Ls=��p�o�jϗ�����?ND5������?5���f�#���XCs ����_���H>�4�<�! �P9Pu��;(��~�XV��y��Zy/T��G6��Us^��N��>O�@$N@�{��u:M�'@�/o�t)V�!��/A]�k��7�q�X`{@����'�SIf�͹\bW<��{+�A��f}���1�6$���
�yb�=0KU:�Ƿ;p��2��P���Vb~����Vo ��(d��y�y{��^�x*��_E�FK^��y�[�ΒT}�r�����@7���D�!�4�1~-�kt��b��`m«h��u�����vSC��'�Ŧ!��y&��!彍�JR�s>�*Ox-����]1�:E
m�D�����N�G���l�����ڲ~�l}ВB)�-˅�7CU�s�U{I7�e�F_�zdht�+���V����4�H86�֟��Qm�f���Q�b��#vu�n��N��Y�3�������ݙ�Z��8� ;Q� �Fnzɀ��B�"�����\t�_|,��Y��%�%*�B�9*�fS��|�'@k��d�[�3�/4�.cOiL*�̘�T8�����L8#Q�*A�ޞ��$�p�5�^�����GH����9�Ό��䋏�o���w�V�����b�R��'��� gʫD�C���[*[���v�VA�-g��YJb[	�P��� � �A�����>��͸�0Q r���+5�crIW0F�+(�r�I�	�uKp!��%��T	iG˝;+p��E|�y��������c�p@Ƿ&.�ln`��e�L�~����*�h��H��)�6-��8W�"b�mk� ���^z�@*f�������2��1�`�*���V��C 6��@�N��>��룚A8��Q�`:�dm=^dnʲ��ሳ���&a���n\p��s�ڞ�M,��w����G+��tT
t��7?<�`8��b�����O;�� ̀�p_2��~In��.l�Qfyw�Yɧ0D�Kxc�c�gt|l�����dcT�W�����S�\��^�W0�C]�@N4��b�\_�Q�Wt	`�ԭ��=y�Cl���G[���f��{
��q��zK{v�n�N�������	SFHLr�g,�5��[���V)�x�'�Bm�wr%3�	cT��x�E�eG�(~�t)�<���>xB��G��!�#n�ϕ�S��!����77�ǐ�T˔�.�Jے"�8O�˄6��F�����\@��'N��I^x�4Y6�AT�@��$�U����my#U�7[��%�Ⱥ[0r����i#\�}U��G�Ia5p���,Q@l����BCbj� NpLC�]	'���(�oyæ	�	Zӳ�n���aD�h@M�Ĺ�Zߡ�f�� �n�^uV$�|�i �=J�\�Q�r$ɣ�U�����s�&1d�k�����]2t6�Q�J�==���z
�Sk].���Uw�kw�ۑ�,����_���,42]�Gd D:Zx�d����+x�ޯ�ǲ�vp*a�m�����gwv�t�`/EOo9��#���f/�C���ϑ��棘��#{�'46�0��U�)!��1-k����>�O3Ex�v�}�P9�o���B���ш�AB_
�H��]=�+U}��y&z�_���y�sn����3#��b�����'RW#�}�Y�u`r%���8�S@��
T�(N�1�ݚ���J�4�]ן$.;gs���S�����s�Y��˝��4��:�&�<7��=.`�0q��Hd��F�Mϭf�PQm�k׹�mc�k��m%
@�����_�@�'gQ��NgT�lK��C\\�A�t{�F�Ɣ����d5��io�Mj�d4Y2���� ���7>*��[�f!��{�p��[�]此�S~ع
cy�&E���4���X�T����Q�ѡ�ȋW�J>��S�{�aDW��-7ut�[��U~�����IO��s��_�W~5=�����zw*p�k��Xѓ�zvT�S�z2��	��^Z�gx<x!��s�L��Ф��vMZ��i��؟S�]�"��X����L:\a����ތF#xl�����q��`���u�O'H��㐚�7tq�;�I3��1zZ���=^��'����.���ٺ�XK^\���f�j]Yؤsw:�|M��=D�ޤQDy�G|��ܯq	���N�q�;뉠�B�)�B�x�����!A�����!���k��Y��!<-�TO8�~����ԧ@�)'�%W��ǉR��(�g}����������lqW�d�^>���ޤ0d�l៘�Hώ�� �0�qE���pE�'b�5��<:�L�J8u|`���Ϫ����"������I�'��w�j���q��25���� ��p����Ah~�B�)x���o�7������}�u��j:��5m[�Ǆ"� �c��I>�K����?T��J\XhC�G��b���F���U�L�"Ah��O4�*�TJ��!8z�Rr�L:���lG�Q�X_�)O�&-ʱ_q�`�
����`{۔��ԼC�-Nx�ҟ��~vK�VG���l��ѓ�8�*@G��vZ�9�l�%�H�)�N�+_���u-�Cצ%�=������w�⏛~ʉ�+)w!A�
�F����u�P+c���ۆtH��R6WH��Ec OG+M�o�����\�ǅ�6b�0DcT�����j�-��2Tۏ��Z�,r ynC�(�E�b�9�L=o��Lp7�+gr	�E�=V2��5�T.�t���i��Ӻ���\�-}����m��t[v@"�(�8ae��	��m�
�N�z?7	C^#�6HU	�b�����u���ހ³���DD�����̔�QA:*$p�W����$��A��H������:W��&�̱�f�`�w���*�|���E��|��	���S߳Q��!�a����oF`c�?D��RWb�f����ǔI;��	�Y No�|bp����c��:��hT�ğg
8��Ù�E��u!�ѫ(��}�ȹ�C�$��>����(��Z�<�)���肗/H@�ޛ#;���k`�op���KyR���L �p��{e�,��7$Sd
���7>�����ۀ?�;���B{$��ub��w��aĵt��i�"`@�EWq�k�ȷ[�T�E׃GOs\X�7*t��W9{jjz��Añ��e��ͥ�s�z�͆���P[��c	�m��r���2�+bڬw��>Q�
�`�|�� \����ùn�cb�}=�i<?�I,ECF����P��s�ָ�88�9&���	����y�-���2���=�$��Ͱ��i�6 g�]������{2���Q�9\v�Q��ue����U�����y�J칹[��-d�U�c��]J;7�3?��j`c����ص��ot�72�Tܹ�%��dq7M҇�u~�##~2k$/��Q[�����ּ P��R0��uZd���E�cs��/P~xgW�p���経�r�Ub����x����=h_S��&��"B�I_Ң�gx�����R��q�z�ݩfv�GO���E�T�r[�.��g���K�{��P2JQ�Deɇ`��ke�tC��k5�5�6�B���,�[�C�K�P�<-��z��U�#�*|����e��[��X�%O��l��y��)t�n���2v����Md(̫�v@�9BA�QɷdlU>�]�e��M0i�^l�|��?tr����sg��6�r��s"]?V����Y���Z����gpƴ1�WW�> \�5��uM 4h�x�R��U#������[o���no`ۜ�q�:~�'OIE�����x��L�a�@yYN�/p/�V���8����װ�&���}0�
�@X�{��xb��&��J�OVS(��#�s�6��<���-��%�U� <Ҫ�mQ�|�H(T��Q��q�-�0���Y}�r����b;`+P	D��.����}�z�";r`?��W��W�6����j�73YM�'Wc�u}YW��W��a����'a*C
�n�S�#����8���Q!�j�e7�!��E�9�9ˢ<Lޡw�U:[qSl��Ӵ�r�tI���L6���N�ղ�s���e7r�>�$8r���ڏ�)��h���w��2�7�0��¶h���%�|0�����a��K�B��9�%��D��J�ЁD�r}ty���̴ƪ���_)��my���%��ܬ�5���H�L��5 ��Ѹ^��D��gL�߭?�˕�zT4�C�%8��s=e�y�"�Lx���lNi7��;�([ǔ�=�L�1r'=��~�s�����ud������kzA:C4��\a�J��b�<@��q�_Mb�Y`��n2����<�ш��/"�.��pfU?�L�{eѺ1\T�i[3Ji��)^����U�������=�zKh	_�pD�-	���j�Q��lK�AY�wNHPw����-m%�(�091��4�	I_���w2�в ~0��`F=���%fY���5Ca�0���d�:s��B�M�Tx�(u���*~ε���j���8�5�.��=�qna���/�}��T��+e�3ޱ�P�ү��s3�op�4D�S�
�����\��g��,�/���_��2��dkJos�؄�Dj����<CC���gz�3 ��l�e9�t|"���MQ��	 ����[�Y/b2�lY8qK`P1�z���)�����ӄ��e�z�%�G�èt��� ��	ޞ��!� }�TX3k��vq�����H��g%>�Y|`�U�C�ex&�>������iTr�/Y� ��V�p�u�O}�*8��^*=�7�+��rc�G�U�$휙ؽx��jR��|��U��ꦥI���ɿ��T�����tm��g	�q�~��IRR��dѥ��h��*����}^/�ڤ��$w�^_��?t!C� �?[2_�P�j{9���k��J��E�S�SD��%<5�9�<�_x��TV�Q&�� ���l�\����)����#�Q��R��<��Y��}�W2�e@�����n˨w�J ��	7riI��U`p'Ѡ��?r�*w�T����񘯛�4c��!�U�Yf��YK�QΚ�%��E�\�����[�P���Ґh�V"@��RCr_�`Eڱ3�t��^�Nn��3�aqq����GO	G��`� �`B���Pв�~�3A��� �����A=+m�]�x���PP���s�ɨ�p����3�CL�jplQ�����y���Ŧ�l
1�(�^hd�3T�O��R+��& ��85}\� %������W�u+�����g�{f��=���N�,�n=���:�e�QT�w�!�K�+�(���/�Lv�J�'�5U��@�Q�9�W��Sp�z��P�/���7����#f���ʧ���"�s�\�#���4�l��>���l��T~�q���^⭨�������u����u�w�.s�`�A���"'4�1�m�E��SR�0�[�d��,��'2�@%�u4M�" blQ�i��Ph%V7 ��}�Ch��I�B��"�;}"�O�ufԒ�*%QU.X���Q=��1���ɰޜ�69���(f�)�O�Л��X�!�I
��	�SY�x==W/�l9�2���|�b��2��2O�y�ʅfcr��0?Ty��#Tt�ă����7.���f�!�O�,�r���cp5%��\�/�`{���L������Z9X�'���w'����ي��zϧP���Q���4/E�%{_�q囕:�%�!��3I���B�Ό���qO:�0rw��UJ�d��c���?���;r�J����9J�W��J�����cxc�.�l��-���4��"�k�ifaݕ�=l(Y��i�e�_d<�N�" u�BkO�����[E��	��Z�l+W "P��ᅵ2ˢ�^ՓEeD�Ym�5��^�&y�1�?$�b�s�C~���To�r�/�G���Im���m�T7��)?X��(��r��N�\P�a{K:��ubp���NL���bZ��KRm���Y9��ZR���[�H�t��z�������H6Q�.�*XudێG:J�"���L�O��MR\�?oj�v�4rf������#4��i�#�_$�F��D��qa!KO���-c_�c` �
��_&�O�4D.�D�j���$������nns>@ǈ�Xr��ULCe��)%���uR�G���m�2�������(|��Ø�T�.���3%#�xD_"�s��6U��9$�'	yz܎G(��D���&\(�����qiU[����;�
V���^��NA���H�f_�}4��kw��C��@~�d��<k1]�u��<�H����}/j#�lD��x�En��4��l������2����C�a�*CxGݱOe
�`N^Ϸ�fg�,N#iBc����̠�He�ař�Sm8jeX�{Z�oU��4v����L�}E�D�d�#�F,�,��&�)�;�{%��|X4k/��}H��Щ��E|Dk7&���Vv3�,�b��ʟl_���?%�<~B.8��(RMuB?]��!K�l�����x<�З�7�
	j���Do�`���5���S\Ƅ ����R�T*r���~1�-�\�q�q�\��T�pXP6>���̒��gLNL�*��W�]�ݷÜ5�8�8u���
�aV7:�t]cX,��5�Q:�+�T5�]P��[�vN%�L����F�׫��`��W���"�>t,}��Ɣ�N����5l֝ٔϲ���oB�k���3�e;\�����ʕ�'�Ѽ�]3�g�]����V�w2��'���������pRϱ<ȃ��U�q���j��L�^��^��{��1�ۨ��ܻM���0��M�"c�����+KP�v�Z[tuNʩJo�xT�3�������fܝ��l-pݑa$-�)�|T��j+@�����:ri�3���aG��	iX�|T��n\��Q�lhx@� &�[��z��7]��������`¢�j�!vaͩ&�f�e_c�p�R%ȸjl\�<R[J�[P?�R�oe2@��S��.YE����p��*\Pd����:L�g��Q+��9�	��A��f�9�����X�^0=8M��	��!�rP�6���z�����g�Rl R�c\{~|7�>�z�jsf�;At����������jU�o�9q�g��d�$gg�績�4�,J�9��igo��w�Q/
�EI�p`��ª�L!�}@Y���-C�<2��_���eFrL�rL�	�]'�8S��D�q5-6۱lR7�G������`q �$� \��c�Ӧ�� ��zq@�gۗ�Q�)�sM7���M�s�Q��g����K:W��&�����*7saO#�-}8�ka�d�)�߫ym(u|�>��,ӯ6{`�;mQѕ���)�}14b�橼7��?�� ��̕���[YAi���`{^�h���=i;�R�]$�બ]����>��f�F�6ݜ����-b
M��\�Qc{z���e��S�mB��#Lapj& L0�䋉6G�����������5찶��Q1/T�r�����R��ʱoZ�������d�w�ײ�K+��q}�c�rw�!�Bjl/�����/�?��ȇ��})�=�&�S^28�Q
���%/@G��-�L����P/�3�@4�ήp&}fY����f�����L�g��>��n~��
��Q�����c��1��3y����T�E�c�_��7А0� D��������B�}%Qc���F3�^"����>;t �P�Pl����ԭ��̻��6�+�s�.�`������c�����D���opȈ��i�P��v�/�?��8�Y�%)�ؚ��W+H�
t�&'������A�=�(�R��I�߁��O�.^	`��N�����Қu�(PS����.���\Y�uD�=�����L���wu�\N+�y��`T��К�'F��D��&ι넩k��k2��ܝ����-2i�*�*
�*zh��*ma�g�nl�1̤�K��f��~���r�*HWvj����J�Ni!�t��UX,f����L;�^E����U��*����r�����60�O��A���e�����"`?�`��X��]�a�}�p]��vF�W�ˤ�;D�Ҏ�L��;�U{��$��N�U�+<�&�����-˒!��s�w�?(����_���g4`�M.�]�~��Y�N�hA~����^	+��b�wՅ�!��n�*EC����-n�,������]~Y��|�`5WU<�cP�
���-R@��t?�2�$�A*�H�Rَ�o���i�e	 �\�(��Ŋ4J����Nc2�"撪Γ3�D�{PT,X�&������Ї=F5D�6����Q��.u'[O�0D���;���V*v*���Z��(��$��Ԭ�aX��t#]�����ںȨ��.��h���qy^�-0�XG#��Ɔ�r�U �2(�Z���v3�r2��1&͔@Ԝ�bW�.t�=`�3�W ��R�.|;F3<��\Y�]��)?�5zp�+�y2�n's��d�eU����TF"/o�)��6'���$����MZ���+���D���,�dw�o�����_���'	�lQ]y��c�KK�?�:j�]�4#?d�}�yc�hW3D.ԈU�K�����N�w "��H<����L�K/��)�,.Dd|tűo��梛�}�u痑���v��Y��C�)����i�d�Gz����w��/������d�� �n��W�@�x�o�a٣�Ak�{3���)W��X����ˀ�z�Lb��A��G1B/�D_���e���?x=	h`jXC���;Y
��Nr7v���)�%���t�]@�L�q�m�/[���.�+��&%Y�6)@	1�[�a�p4���Q̄��U��MAR�u�h���pF��Æ�1��(��ͅ�}b�"5�xd	�hs����3���.i����lf���]��"�?��lᄃ���Gu�N)��'N�d�ت�l��#��y��w�]DC_�_ǟϟx�`�VcI�v�h��<���j;�n���r5�G�Y�c�F�mO��ж�s�+���>�,�O�jz�68�Th��.U�@8ͥ�����vFt.�@\��c��O/�����h_a��=�'Z��ʬ�����%�(��j�`��l�5�g�9��>=_�^6�7�'�s��#Ny�2s��ehZ!��`���_�L�|��BwP��S�����Y�@�.�}"�����I�-#�@�t/���:�N����6�k1�I�1���P..�6�OzE-��h(�&���_a�6��5,U]�'F#c�c�y���]�D��~��ɍ�T��騔�"4��=ͣy�QE�]��`�,�%��n�u���'X���v^󃍩�,�3U����h@Yמ�P*����p!)�/�2��;��"�E
ãd��!]1�߳�I0���^b�&:�i �W�p_d5{_�����쾸RWm=?��\�����*�U$j7Y�7u=|ZF^ɖ�f�F�q<�����M�܎�`����Cb>aB��7#�H��q.�0���ʌ\�nr��I`9L�	P����-�Ź]�>v�����恐'�PC�ؠS���b�9��
%lˠ|�(F������^9�Q��&Οd����J�����X���p� lJ���b8A�^����>�	Zx����D$kb$�K��������A�cw{\��bq��X�g�������ĆA'�xZ�oY�͹�cJI�t[�K�tT���A�j�@��/��yv�x�ۂ�-�;��� �.��k����/�nn�%�Փ�0�~��y�K�;��J9���ސ����8�A��Ҭ�{4u����p�`v�Xs��ʲᒲQR�n;#�z-�ÓU#v*��q�n�I�%jJ���c��n��V;����7!b
փ�N��ĀKYA+ݐ�������X3��3:����p���vT[�S��v�I����Α�=����j�|ĝ�V\�WR]h��?��1[���<�g���h& �Ƴ�x&��񊻨R�
�����We>�ϬV�>�I�t�L/�5�EӁƠ}Ρ0hlq�� �v��4��'��#�S�M_ӧ_<*?�w��3�� 6q3���D��WW�gOM	����[!��?CaN?Q|����<��@�F1�ZBX���J��v;�����<�9j<pqH�5�=`H��xA7��Z�0c��)�euU���vHF-0~h���g:���f��d=2�"ʁyŒ^/�u��KRU_:�&=��`i�A��ݪ;S2;׏�j�i�RT�<��z�t��ԋ�d���hlX;�$���>*+�öј1��|����A�ƕ�kތ>�-����2PG0��(Ϊ$ZtB����ÛC����u8��9񼱇¤����UmY�[5�w�DQ��{��*���S6Q�T�wS\1!/ƞ=��cs�Ij��k���?����m��Y��Fv����˼4o�c�%X4��\P%��I��[�+��S��k4?[@&0Yyv�OǊ��7�d ��Z�EjAs�"��H����wW�mk8s�G��-9	����'\s��_��@o�2���7&����Oi�h��'�{�c����Ҙ�,���!��,ٶXX��߁m�.���[�yY=��@�
(�ps�|YG똦���־];�f�ZU�b�y��h�j�M�����zMt��M١����	�"�D�"x�'�P]&c%S��� �&��r�3�g�x|Y�J��ʱ�kĈ��;�琨pc��=X�m h[̮ntu��7�	 �k��Ĝ���)P�� �с�0�ښ�_��}˞:�3N��Ӡ�`α6���	\ϕ�Y��-��m� �tcW��+wL
��x�l>OljB�
�Z��.	�o8
ք]�T���I�
���]�}�9DF�rw���^�p��c�L�ϧ��d|��_�vĳ�G���yZ $P�����á��B�x�TEk�q��u��T������x-�Q�k��ؚ�wڐ&�����isrU3�0�<�{&�ѫ鰊t.O���ST���*�� ��N�/��W�13���`(�*�M؟L�����+�)�۪��
FQ�٥�'ڪL�Gu.��
�)�
��iۯ�C4z�j��g9�ZY��s6R��޾�4�AjT�՚g��!��m4[��5�I�<���Hc�y7��X?(����}3�nC��3�Qg����wmka$
d����T�G��<9M#�!/���ӓ�V�������|RV�����Ϣ
i5���Β�xG=����W�ij���^g"9�Ă �����s&&Za�7��)������ٲ��@�-��Y�"��C��k
MM-z�����;��>Rs�<F���m3�i����*\�M�>1��W�[D�%�onr�f8Z͡rv�[{�������� ~s��p��
�m�3ܵ���>=z�v<1E�k��Zx]#�؛/�*,ւ���@�&��rѳ��ԠG{��z��aT_G	��4�)nRY���e�2�Lǆ���쳯'�EޥV�k�^����~�P%��70\���M�h��<^�"/wNј%0�$��d#+��"�^ ˯��>ʝ�����]�R;�|��^ŏ'[��8�L�S��֕�Rj�Z��>�HH���c�n�!/�	���\����*R�!�`�U��2M�r�=�2e[l$r���ӱOdJ�D悔��u�PX����k=k�=S=f�	���t����~9�FHhK]���z�P��W�Ʌ��|_�`���́���>j���ֱ�)o����U!��W�1��`�*�k5�������R}>x�޲+=��}�70_4�<���Kz�s �h��"�~V��j��(��R�ȴ���T����r�
�=�>G�M�>�|^Jڠ����\�.�D]@�aƘ�I/��*�'{�]��G�(�ݙ�-Em��:݃�4���68akb ;�&�m4/�6��yz�;�<T�J}�ա�hKN�+��x���%�3��=A�z[� ����i��`Gg&�\���#�|��W`~�x�nz�����s{��"V�r�O~O���
�`��aR�vD����b���o�}I<�ؔ�V��C�u�6,�toޘ��� HnB��\�U �n�o	wt@⹬��*��1�7l!��G:�S�>$Ԍc�XR,JG��ʓ��X7�+����,�m�;�~�gs�c��rt�F���t�'�U"��Xls	&Q*&*r�[&,�}JK�ނ��kJC`���P��i�<����Rd���Q���C�]&`m�G#�)��tN��v�(�c�죙�����:�3Ԝؑ4��,����a�I�BI�صPX���מ*��z\�^��n�L|T�{�e��~����E�V�.���+1�S��+gy8����ё|�����<��Y�@]����Nɻ�:���	�~ �aZ,%�0M�鋾���̮u0)�)�|��^�7�׬rQ�X|	���p��R���]���u�!��{��H.n�Q���mnBD�a��v�j�M�y�ɠT'Vu@A��ԢyP2 ���;����L���
��5��k^�
������/kdDG;S*�	ߠ@l�R�#K��Xl%P>%]!�`h�4B�1����*�_�|�37��w��Ƽ�[F
�R���^�of�L��;s�1`<R�3L���!"�?�0�9g�����M�N�Mȣ>~���2_k�7��_Rw9f=�lN���B�kgw��$�;+��NxޤR���LG�h�Nˮ��t=�̎)�w�M(���̭��k_����WbU�ur���	|їH���3XlQ�c�� ��.�ihHa>�����s{��s;�d�RJ����پ꼣�=(2�O�����&��T\o�FH�YCj5�JP����Ԇt�8��q.WJM~��h#߻3τ�i#�I'r�J�����s��l�#�@ݎ1�u�("&)r.\JY�Z����g�݌���Pm�N�4W�U[l��y�55��"��]�fT�7�{���S���5��2
Y	N�����p����
����9S7ۜ%����T|�𱆬b��'����>}cǩ�Yꙕk� �G\قg�����ٜ�#gA����*<��&1T��.�t@Hs���-囝�Eԡ���Wl@(
�N��;SQQ��-Bbd�e��`
�f����������OR�ۖ؎�|��;��nI�������U�f1��S�ĝ����鸎���D�NKs�A(���}���T�+�z�:0\W�Ǭ��HE}>��~�G�VU.Qsc"3�U�y���4�bs.<���.�Ĕq�_�N�U5C������9�4�"����&]�7�a�����>m��l�cd�d`!�+����Ii~�B(J�)�L��w-H�$�IF։R��#\q�e���,����o�t�0{���'mB3��t�;�&��X����~��L�P�����F<���ס��4	�4^[|4�~J��Xg�`�ٛ�&�fԁ�Do��wP�
���ãa^�^2û4�o������.ힱ��-<��G���H-��&ە ��k�����&�����޼�M�Vb=�8�'؁&&j�3�z�Nw���Dl��sf��P��O"I���v����������3ml���(��]�)DH��lJ��g)Z h�!�W���Ճ��A+.��/���j,�b �o���i����-�r��p���;�g�0L/�N`��Y�w�t&;ܑ_��i2�Rbk{l1�f��a	��.��˵�$����	elͶ���D��+����+,\��VX����u�݄LNuF˛�Z_�J�-V����Q��R�ׇ��\=\9�J��wh�#D�.��>9b� 
��a�����d����/����z7���n���A_Z8�$�R�s9]�(��[���h�pX�2p����|�on[ݑ�%���KA�)9����݁`⮚�5M���(��[�|�Gl��~{(�"��p}bEm<�M�J!�9���Ţ1Y�M�Dc��j�IB���9�v�����ϧ�P�A2j�u:#�\�8/]��޲�*d�a�b���y����EI���< ��.���W%��m�w��ꋌ�`�%vAtI��Zl�4r��$Ν<�o�qg�'���a�E�j�4���m�C�~�C6���9s�(�Ѵ؄�Z���:\�>U}��c���YDB:ʓ9��K1�2d���.�����l���*� 5]LW�ƢeqI�|��}weT�UVO����M������&s||��b��1{����-z��J��j���,-�m��+Ǘ!�5�����rI�K�*�o�R5E�P��3��.)��2#Y@Tj��t^�_�	^����� q���'iC-���F4�X&���?�L�n�h.�yO�`W��g�c�f
��g(��g�lZ�u��R�S���,�'|�ʰ
��m9��������5�-w�=�W#{�N�.rڪ?�aq1���MQ���v�G9��9����.��% ��^����G������I�b������Ǵ`OѺ�T7�k���5%E�������m�}�0X�>J�~�"��	O�������Tǁce�����3�l� T��(w��^uє�p��|��k*Kx�L�m��Dp߿�}�͒��W�:�8�3ÝgsM�����{^B
� �n�H�U�7�/���#)p�n�xe#�p���tQ࠮�]T`�|�xoi�i���Ž�>q�R��H)��]���.�bN'}�.[s90���X/�`$λ��kB�N��/��:*��(�	�~�C��x�,w�a3S�^V{7�/"��ג�R��g�aPBR�	j�d�_�rz�k##{�/�*/����W��7��&R��'��uD�s�g���gS��rQ��_bI����c��@��kTp�v��ZV>��2
��������B�'Ǽ-�s"�Q�L׏��Z���%2r���V��ai�N� 5�Y�+�52���[�f���:Vd �&�wc��;I�j����O=\'H/n]k�P�w#��S���ͱN�R٪b�@��ރ~5����V����&RW�������R��@�� Y8�lj_	���H�R'��熡fk�H*=���&OV�p��k��D1�t�~��������O�M���#[�7a&	B�GQ��֨vT�A�ɢ���n��b��� �W,G|I3E�2���C"+̓�)z)+92rZ(��[��Դ��2Xw�ĭ�:L����a�9������+Fi��k�AL�P��p|8!_����.�ў��Pe�<57O����ON������S]ζw�=�'�o�!�\�D���[	\#��#���U/���2�N[��y>���&q�T�)Vf��֝F�r�A�ٷvZ��Cw�ZtYrj�0ȟ�N��;���d�����9�I |@Z��[ԏ�&xVխ))�}�.V��%�� �V'z�55P�	�ƣG[;U�9k�����ױ>wB�ߤOn�R��>�,=��=�%"]��7�=W��?��x��D�i�"'��ߍ�5���s��*�9_1U�L���r(�ʫq�5��'�U�,^�ƅ��<NL�o���О���!?����v��f5� �g����zu�����λRg�L���=�UN�38}�g�3j��`+�Y��p��!p&����T�d>M8���QЈX����HBq�t�-��sL(�i�Ex_��U��j���n���ndZ���U���c)���~��Z��Q$��Mi��CD4kb�������׼�NU���5��J��o�_��Ӵ���MQ�oy_��U&��K�cF��(���JZ���v���1��]��C"�y}7.�>U��ڝ�aj |�	���A��I�2�q�' �w�$E�{�]�(����?�y{h�M3�ᘓ�B���zªA�_������yL�[��;��T��$3����/�8%��������J��2.��Kg�zp�q� �Z&B�ə���f+C����V%y6�jr������"���Å����·�C��?�J�f�c�^x�[`�m����~M�����~3�o�K�~� D̄;hq����
ړ���PW~P��ˌ|�7��aw啬�:��L�y��`�i��*)��Ќ5�t��֏9눾B�mjy�}��O��:��FP�q�a�&�{��3���t|yW�nE�qSS��.7�G�8��G�t��2��4��Fl?$CY�ȫ�*C�:k�Ԗ6(Sg4��腿����2:ɴ�G�!$,�A�­c�����Il�3�h��ϫ|�S�9�h�����M�����<��	���h1��f�O=�t��ش!Ms�d��B	�/Åx�>�T^n�Ts��b�歝��"@�	�mq3ꕴ�LG��p�z£��o��B6��"����W�V;�FF/~��A���*�*;�ϗ�<�#��~��=���/&��ˠ���#��a���v�%G��8L�8fx킋=)Pg���Q|�[仾�d��T���򦢎X��;2��C��J&c�F,&ȴ�L�#LV�s1�j�k���l-v�f�3���R�#`\�gע����P<�TBK�a�UKc�`���@@Q"�X��@�<�ڛ��:�Xɟ�xR>�Mdի��&��� �$w�������4����Ԯ?>!l��r��M�G�P1�]��b�j�6:* x�2]:��ٚ�^?�:S���0�Hwi�\��x�Ɖ���x��Ee�M!��]-���O}���uVWqi�\��&���LWV����"64\��>$�Ē�.¡KS_��T�C)џ����ɴ׵^��\e�1?���^��ֹF��|�Q�����!���$�w���jQ�e�%Y�L���e)�������%F�^ժ�2�5H^d@�� �{!S:�W;���&Л5>˽�
-�4�>o�&�2S(��Nq"_�Ҿ��\K�Qm`@�͐^���HF(���Fy��0o��<�ڏE*�r!�����{)9��m���	0��S���*�I�'�h�FCb�#�A�MI�Tת����g]Ԛ�XH���=��x2�92�cˮJ�cˣ(�Qg�)KǼHy�@A��v�����D9_�:��Fe��m�~(jNMveƚ��lY3֠���_pmv���?0�c�e�Lor���t-?xhx����8�S��ILf���/�Ys��>�rC��8�k�KH5t饍���������RN�=���z� ���Z�9��#
�c�w-�Ǫ7�=*��s��!�$s�6Q���0Q���Ԩ{�c�>V;�ְ߯���w�y�W�db"!x�hh�>#���m֠�Q����eiȹ���SkAZ��A�K���]��2�튽p�6� ����"=���r_Q�땯�2�^8J|�;��$\�^������Y}���Sb�m왐�n� j��&��LC��6������l"P�,+B����a�����L�Xk�)�E��mw:Ș���N�qd��*~H0�oB�*�l�g���m+zϝ�f8�6�k��|��Zu\��P�d��GwN[\�z��(<��`�����]���
E�D괹4��z�ڲ�� Y�.�������D֛�k� sQ�Na��n��{�e��Yn���~9Q���h���Q����$ٱ&$W��k�H?]��o���j�����zh'n5W�����i�!��~r�B��(����?L�ќ��L��(٧B&���h�p�U�ZV�!Z��jy�˴W�-=�H�q�*B�fD����+��8�R0�O5�n�=��J_�%������g�82�A���Aj�N����R��Ќ��[h3�{)s֦�/P�hX9��7�=0�21��De����"����D/���pޤ1\W��gO�hk�(���'D��z�*#@�3z��M�?���P#�)���)�8��M=7����Jk"5��9��/t�U��O��O֖��b8.�d:"ӿ����v�h�@"HyK��B|x5#'�a	�E/5a����'WWSے^	8q�@���y���|��Ð9���"�H��Kiɵ{��"�'�Ak�Y��ט��븱�d ��3����AM�{�eX�#qH*�!�%*�	�`�w�������Z�����]�u�M�m��[�!�����ø�}yn]���-7 �֋��?o��'o3���T���Sȅ�dT~�>w�fڹM�+*NW�O���؄�-4h(�yjƌf JP{L�I�M\�+F3�$ik��]J#�����Q��x蜉}Sogp=����{�d̳k�m��+�!G���Ej� �<Zު����u��3���_L�?!����,�$)EX��/̐�?�9�˰A?�@f#R��_�}|�7�H�c�������Q�t�[>X�f��-(6O
+��MϹRE�5V��)l2�W�xL�z<��5\{6�*�-���&�'O��_�y�I���aP����9��A���i��3ْ@�����@�Fq�V4=`�]Tl���]xW�,���l4b0�c-K�YK���إ7$��$$�xL^e6<�=�ؾl�'G�C���K����S����v��5�E��_�����iIl�mX���_�s,�>x�j�-�ܢ.��@���3gC/#A� F?��dm�v���J[����}�Y: �fKKsܗ!O��z�ɾў:v$��$l�6?y%#�Lږ�poa��U�'��1��'�:RM���9q�jM�@DK�������aѮ?>�`י�o��P*�5�w��n1Ŕ��Z�˹k]e]�^U4��S.�$�/Amu��G�5g� �HR���[B�j���u4.I����n�|�
������Eie�P$���qd�G��k1�Z�g7�(0)k��2G�Hx�ٷ��Ol��Qz�u��f�P쒸^�y�D��'�skj�*�툆�>��_�f<?$�]��\�
�&6��!��[��2Ĺ"蒆#�1y/�Ay=Y������Pt�/8(�(%�1Yu$娩���R�!2`C�&a�H��DE��}�z�x�Rj(T!׿�7W���Ȁ>gPBQ�|��������hb^{��P��{}6l��|~��=VG��n>ː�BxO����o��{��5Ub gL�|�?<Ffw�y�'�S�~�����j�������F�1����#R>����R��� C���Z ((M&��*������V�\�;ք��=m�۳4΁�,"n�-�w�i�`�� �M�\H�x��|Xi����UC-��� �����n�n�]�KC�w���"ՖW�	�>dGQPf������K?FCdӨ��J5	b	�C�ܑ�H^jQ��GKP�L��hp��3���,b������[��2�/?�\���&Bj �]�/آ�ݧ����aR���åC���>/vA��`b�
Cـ��o&7����St4�ʋ�j+[3�K#m���7Zx�mrn!+6E;Z�ж[lH|�M�o�T��j��V�n1Poy�[�1��}O޶��1�,�>wYMe	�b�ۏ6��5���5�8 }w���{Zs�]v�Sp����XxJ$�����.N�� ��?���?���1c�6���g��ݨ��&0i�f\�ED;h�PN��V����wV��8H��;�q����V�〫�M"_pz|J�����{?[��7��Q�k��gDB4M�:i�,�wOk��̢�_y��)V�0שD��Y$�ԃ�I�?-�09w��ҁ�Z_%" ���v��X�Ⱥ��
e�x�
N�8hq^;d�F(ɞ���+f�G3+�S�o��J��~x��nd�\E�7�W<\i��'�.$]�A�dA.�I���ʜy�ѵTڴMW9Wӊ�!h�f�3X=���+2���<Ȱ�(G�C�7���Վ�7�Q�0P�{;�2y�����L͡����q�L�K��X�a�#&��^Tlw 왼*��ײv�����z|��C��؝�Ӗ���m^L�K�`q��_ŉe`��v�#��Cp�������)�r[D�B���02�w
�,��hG(� EC�-�4���B���K@�ј]P�.e���C�x�-�b��#_��V��ő7Ў�f��U;��c�������!����.�Ei�<���
��(J������L��������~ǖ&���.�Y�˶�O~a�+��U�;�ԟ�lp�dM%<��||�s>�ڱ>����rǇ�2�&�sa1�אziB�`G����)j�\���l���MZzY�n�#�;ew�h�8V��\�͚%��q�/�t�b��lZ5]��:ym��|��r5�2��I+����Sn��U��Y���if}Vz��/��PB"Q�*��$��&>^�DG��<�JZ�����tԃѷ�Y]�CF����h�Qto*�%��y>����!���2�9S��i~�$:P~c=r��*$|�G:�'J��K"���|�|Kt�^�AO=��Lҳ��?�������Q����X��"���bs�\B"ڪ�X?z��9	�ڥ���
F#����<��2�f��b�3�Z����m���Z��g<3ɒUL�σl��DY����؝�:��X��b�g�k#��R�?E/�jwN�B��y/�J���Ñ��|�<��I�&��}Y\C� �G�{A	/�dҝVU;e�N:��#��*C@at�%�(m'g�ֵ-ot�7+�v�S�>M�_a��+y�ܝ&�)tGsx��OQ��Z(�4M��n����2�G�����D�M��+����gSf��B+  7m��c4R��8����f+�u���-Y��1��j���((�ьM��P"�X��� a�~��2��������.k	�]1��2�āU'�������UM�T��4����o����#y��mG�x��d�[�>�l�;m�:��9MlRֵ��Q��y�v���N*jg�^^�;A�I0�A���!u!�;7�9���L�F ���ؚ�4#�ӓ��:���4� ٞ���c���l��Չ�[X�]/�y)>]���e�jD�D���c����so���,M�j\������nym�����n���lr�6�,)�@��������CDg�!l[4�i���Ew���t�>A*��{�������y���uJ���P����\�y>��?���켋������|�s�0��>�3�;�W�jǴ�;��׻md |% ��<��Y޺�"��:�t32���Z~%
؟*�j���T�*������a����nD��_��}v�ȉ"�o���ZC6s7Q�6Wq}ų �W^�4��*TC�0wE��L���i �=R�y���՛��Zq���H�m�ʏ�1y#1x��q�E�+
�B!?����{��������}~��JF
��� שǓl���p�3����c"8l��W�?�+�c���!ϓYĹ6{ցi3#��b�l��,B/p�e�n��֩]gD��ؐb]1H�bI�a*�= D����ev`��Kd�O#�y,�K(��nfy�ؐ��q�'Ms���}���l)>P(b��bD�i�,и�&��n$�͙^�_� f+vN�Kz{_t�
/kk� Ñ9x�?��n�v�QCF>e6�y��G������;��=�,�=�h��ћ�"2A�(d�����Fe�c�Ƙʮxۙ�;}�ܳ.?i���&C/لoh��yLr�U�ǡ"<w$eԩh��-��]��By�D����r�isb:{�������+[�VQ�Avd31o�5q���8F�s����Ӌ��7y6e�s)����|T/#���,P�U�����~dԒS���[�21���deP)�=�j}R�+������X�
���j*�=8EՊ��
↹oT�G �#�"-H{���(��� ���f���%/(�B!�Eɜ�.}���(��Ñ��}=�,�X�!?��Y����%��ܟ������a,�3. �K���H3�LԪ�C-�ٖI�]GB.fט�u�v���D����h&^%2S(%^���
�K�H��OK�d����§�!N�p&wS��z'�+���2�w���ӨZ{� C]o-q��FvW}��ٖG�d~��uW�~�Pe�\<bQ�{5�Y�1 ��m@]�E��$ľ�ȗK��g��73�X��tS/vK��Ɲe������op���r�$�xǅ�'���;=LX��j��Ac����B����O�x��H�~=אB����|owL�=����G��f�>�<u �F�I�fQ[7��9;p��$��b - K'����7��ٿ(�������_q���5P�S�6'Jn��T���ݧJ�#��*��8�i��#B:���;�v�ښݕgz3@3mJ#>��H��e%NcN{�:���7�Ւ�,}�ֱZP�p'��J' [��� ��|�'��B�_
��s�9;�:sL皩S�5'�,y���g�O������U,�1��� N�Ec4�9�I$ѭ�o�5�Z4�����||��B�a��D��sZ<�_}1���#=��-�P]ӊV�z<�/'�q�[tC��I���o��(ܗu.lx������2�b��w�C{p-���8���T�^��%Nn٠��L��Qm��־N�T����'%�3e�Y�Z����W{H�G�a���'�����X���|���S.�$��5�EM`�T�Q�D���{���
H�K�mfK�wЁ���΀�ͪ��ܳ���!ݧ���v֔�K=��֕<�/�1��ª^T�a��#շ#�D��w�����-��m��b�t:���a�U��r��cީ¾@�ۏ��-ڜ��l~���7���HqN��wI��ѣ��2�i�@8���ϖƉ� �+ܤ&�|Vh�f̄01��-ާ���L�o��U/�����݊�B���J�ꉫ�(��)V�9�X�o�2$���zU��{�tc8<o�G�cgQ�P��q-W|*�Q�|3��iH. ,/��7����o'�0eʃ,tV���)nI~���H%�R�܌Yˍ	
q��Fp�8�j���ݘ����Y���Ҙ�Y9�u=�󢤍'.�CɊ4�:3������!�b�u�C�-|�R8�|E?�0� �,�V��3�8 �������~��q�~_l��X,�zF֑���k�����3z&xQ���g<}�K��t#b�Ã����)u��lK�D�.��"m}ݓF�Y}��B�C���ww��z�iҜ��f���q�y%D�Q-�K��c=�2 $����zS��,a
ܙI�E�Y��k���8����O����y%���m����������-Qĥ�	dc�{UO�jQU�ߨ��K̖I]�t%��d�������D�yq&�Jw'FM���X��ޏT Цg	n�5������r	2�^zT�]����ləu���m��D�A��81v��[���Bw�PpG��m��+������p�12Ջմ5�7���nww$�S4�Uc1��'�l���
Zq;��:�|Xg&�ODA$��T%=!$4�i{؇�����'�O*�Ѭ��rkq#�b#ea�"=�7��@��Fk��J������Ң��&B	�5VRh��lc���yJ���g��l���c�ف�	�(�lӂ�Kk���f���L����U��.��[a���|Y`^���*�CX�#�z���.�k�TZ�A�����e����<�1�#斸 ���샿��(Ysv����#�����y�@k8��$�(�.�7���݈Ɯ%(�%Ww08��LiU��W��T v3q�Fq*�xQ��+ʈ8ȧ͋��H�m�"9��m�y��z��~�E-QV��ʫ�.�ٍmc�)���
�����Q��ckT����E�f�h��7����,���-Q���C��߁�ha�W)>f�F�Ԭ!����#X�4����YR�(��E�"��z�������?)���<m�+�9��сl-몀�t>��չjM�^L讦P^���(��w������P��Xv;H�j=��~����4��E?��<s�E��4|֙]�M�<�B���'(ƮcBu���J�;�|��<ĥ������4�.�P�hZ|V:j����&�ݸ_�1���^G~����9�5����̜�0��a�<Y����v����_�`oWHX���<i I�T���9i��iq�'�.�=������L2�|�L�3���5�[�8�tE��o�=�M\��L���#�D�o�M�\BV�z&��5-t�S�qI��6����i΀B��9t"����X�S�&���0�B������F��s��gpt=���~�F�_E\Tdn���<D�F�1��� �B��J�C"]������f����8�K�=�d�&��&�(Ҥ/�~���=g6��f�wiq�V6�=�	��p&�� �Fs1���AC��DPzWze��� ���*TQ�n�h�����$=]<�a��т��TŖnR�`G��i�L�Un�!�Z�O���G^�v7� Q�T(�*ʲ��+�d���1�5�g�
ze��eȶe�^���o\ܺyw�^GL,�"���a�h�HltW�Q�ɟW-����[Ks���������H�����3��-':͏��i������S��G�V�K��x2�uGL�L����]Tf5u%'�@@q�*��v3�K�6�oL[Գ����x���ZQ�r1��cz3�r���T�ܞac��f6���7V�g
F-���  *�)e�|d[`H�1�B��.���90��q�"�A�w̛�{� ��؍?Z�-����n/U/��O��.�Z����kN�op	l#ɠR_*c�B�R���=d%�Qj�q~(U/��+��/&���Ӻ~�o��˓��=���\�� B�P��)θ������ZL#�v�33�7��h�~��5����q�<:w�q �� f��|-����"�HwXxDE��9`�d�>��J��m�0�r	���.�������h�x?�9G)k hJ��*���8��R����KfX�^i�=�胐qS
eB^&}�]r�wl����]�5bO�.���j�����]�4���>�8e#�֤�Ev��w@���ߚ�^=������C��O+��f9�nMj>�$�����(���|�$,WSn�����1,�vY�_�� ��X4�g����'_� nK�֢�C
�b�J�5��D�ysE,z�����,�N��d��)x�>cS�P��Ӳ��l���M���J=���'���lӥu���)��_,��#���U�y�?�'�ydX
���4	��i>��$'�)'ER��>�B�іУ�iW��k��F3����z�X�K���ۉKK�`OVg##�|Y:�r�5�����$e%j)��RF��B��R�ux��e�Q�D2�(e=��^�}��Z��/c�G��$�!�t�o��9|���-�KãPǧ�o�L߁&Rm�PR��T�i`7}H��KO���`5��lLq `,ɐ���^�IVP'9�8���h����Q�V����t���5Fwg�r| ��A�j)�����,�d�W�v֮�0��j�FV�|��a�l�)EQ`
\;%c�G>\��������X��w��.�v��1�8��i\�r�0M��+Y`H�ɍU�Y؜0 ���8@�2V]vޕ�__�ʱ�28g�m؞�u-|�;>�Tv3���(�W@�@�إ\~���CC��o����aϚk�@�A�Z>d�7r�y	�h��Y��<h�c����� ���:�	md��M�Jp��|�64B�ޠ.���3
��"���A������z�z�h0Q�e"v&y ��,�P�ȜU�dQQ�`E���~o��P0�5ۦz���(�d4�[���o�_�.��ܒ��B<]>Ie��WXv�R�'�������&��G��	��CU�8b��M�C
[;!R�ez�|k4��(�eX�ë� ��N��S�陈ݹ�{�����K3Z��y^�Q쳖���Xq�Պow����5��:� D��NJ������W�׽�����j��E�-��<���z���] ��x���F{e�&�����6N9���R v�����N�����l��q���V�j�JYe27}����)����-;%{=i�����5Q�m6$į�nb�oG��yٙ�՞�
3������t�j�s|�����k��R>���Z�$�b��O�[�=u���}�A�Ǫ+Z ZK���~Eʫھ���w�v��]C�c&ji%G�S1�IY5q�ǾB\�pI�����筘��:����!��@�l�4D1g���?�uT��ߖ|��OyH��M�����Пݲ��Ե�4fo�}N�Q��ɣM{agT� �5���dY���N�V�fRD�rGvd.���|/i>{��)�O���RE���X���yğ�7+��>��].U��C�)3�����_ߊ��ˇ5�x�<ᨢ�4�U}��֣+�_g��_��H�e�O6tc}V�b���˝s��0�݈���[�)�_<����Q��VmǛv#�Oѿ�B�co�]�n}��6b�������ԟ�N��Q%IT#�T����V���k� b��3��`�,�XYQH�$��e���{�e�<�3���銜�.�������Z�Sl+�՜�|��\d]i~�&a! q�>��U1�(�6� �]g����5�������J�c!&� ���������h���Zh��A84��O���s���}:Ø�k9�Ԥy���k����V[���	O0}�j�JV�(���{���u��3��nT�qî�l�������fa	���� �]��'�QD�y~5�{��^�W�����"����tn���J�P;�h�ǓX2X�/�@�va4m���Z\�߮p۽�[AOf����[ +���+=^=p��P�&��Q�k�����*E۷��2�4M�Τ�W9F���S�6֨�E�bv��ň�OR)�TH��fFJ)X>w+?i�<���3I��2���.��$����.7��	��0r�ߎ�p5~�� ������f�i"��P��b%!*��L���O��;� ��S<�=�+6�����}�Ɨv�B����fҧ6uPl�|��C0�Ϛ��`�-U�澹}�ߐ�Y�+6@$&'s�-� X �7�j:G��8gfEP�'f:{Q�@��������f�Y��w�mZ�(��E���VMx�U�-7���p�0�IAl:l)A���&a�'���YO^��"�T�:G�cfr�?��`��Ǔƾ�'n��w�HlW�P�ɾ��@������M5��m !�p�-��1�$9ElB���XWG��9���+!�4J�diD��=�XP����W��|h�a�i�[^V:���"Jl�v7~��c�̚�F�bS�"&��5#0�(P�[���f1�DG)�F4����8���O�l�V�~��L	G��ΜX��Jj���R0�d�i��頻�=?�I)����1o+�Aݟ�M�/%�Aߛ�WD?2G���F.�����L�ë��'굛T���c]�PX�;�@m/��)���9�Z�����-�ĕ���x����J:l�a`.�����?+��l���x��{ez��骏�a�(��A}s�^7��2Znu��B��5Oh�"�؎W����p�+�>{�5¼�/��)><n�%���L�j{w�q/+���ŀ��w8�nw��Y�u��\��,��]Π�)���v��jcp�#���#Ic�Ʃ�u$�O7�Z6��0� N-����61��n�N�I����e�<KD�+9U�fc (%���'�ɏa,����v��5�'���x���x�i�a� %ph"�����d�
m����6���w�M&tG�w J�ϔ��%��V_�l���ԓ&`��ܹ�"��Bǻ�f�-�.��e c�e���D`%���@Ξ=#�3���_6�NUy;��=&{,����"� !>6���/�	u��x���i2�
K�s_X\u�n�|]c�q&%����m�b��Л��%#AIw�[�\���Z���k�?x[4m��Ej�g��O��-C�"-׎h���SƹRi��i��W�����R����O���ԷS �YP�b��ҌA�_ K6��v�y��!g�Q����
P(!*��h�Ӫ��'�Α-�**A�9&�E�m�U�y1R6��3��ğGfj��y�����h]5
��Ҥlc��1dr:fXj�Z��4S9��jW�SS��>Yݽ'� �w n-w#æc�`6s�5���&b�c�Pd���
b���i�׎��Ue��r�@���˜U<�c���e�31�I�e\&Q *�!��J̈7O�5N�g���96��T����ft��m_��^GM�pmT�?�vUBe�	�n :�vc(-���y`�W �ͲG�C��gx����b
&s�S��#�D����%ׇ��-~��k^{l|�dA?�=% �j;�:�FKB�H�ib�7�9h�����a�B!�dX�Kg��4�a������B�"��F�~w �:O8`&����tV''�d�)���L������RTR��Z�S	��d���_,(W�5�+o�8]1j*�H^10��d��.��-"қp�;����y� �T����>YL/
Q�)4z�.@M�ί��67�#� �PvB�j隂X\Mv�f��H�{s��}nXW[�7)��`Җ�$]����&IG{ža����Z���\G���
9�3h"XnJ����ts�*t��T��~^`m��Jy��,���u8�WT�D�Kl��>z��C�Knz����M���ALؘ�YA�:Y���A�j���o�(�B�o�u�0.�c�-�J)m=��F�bZЧ7�E'\�;f�/�^}+;-���M�싡W$PΣ!90k���{�t�98/ȏf�ȇx8%�~��S��۹v�?���](������˚AZ/�X[;�B2l:���L�_[sվ�F�:e�8##��ĥZyS[���w�e'b�� �ɝZ��;V�J��g`�`�����5�Q��ȃ*����\"�H�f�q��fR(���J�^>j�5�m�E�"�������cc��C�u�n*Lwf�+Al��5qʳ��4(l$���][h��#���3���7k���p�u�:�m��;�]����e����r��N#!���u[������A�]� ɦ@��Ӎ �y���j�yr�[�XǫQL�� )(��c��	t���rs�X{زi���-Qq�2v ):��t+0�W�o��<`@Tk|�P�ȼ�m��̇�T.7�%�!?z�{9�Q�ƨd�a>�a$�t���x��kS� P��Vc^�A8Na7���t��>>���r��f�.�ێV�|.��}{��xD�3f�%0g�T_80֊�J1�5�!����0Z���r�y�*�M>J���6>���:���d�i	2�K
��KG�=��T��P�m�*�=��˦ ��mcc��_��0�j��}�u��<"9��EU����T_a���;�8K���0.� �빲�4e�e.������$�>�AW�Zr"A��i��o���7�,�QA�|>-��9���!8�0g�K��3�lo�6C*��K���f��[{$!�À��*a\ޑ�N����S=��>J��?`³o�E��~��y�>��r�)H+�Ҁ�B����<0�D�&e�H��y-*N��n�'�%�.�e��`�/�R� @ai��Ipp"�(�� �����[��Hv,r����Y��������$�{���;nV5�+r�@�l��ՠ�d�r���}��q���kL��wo
[����z ���pMa�v���B��]�}�$��-�[���û�%����$Zj� c��7��A��lP�Հ8�Id
�U�^���� �<M�f} ��\���HW��j��F�Z:3�3>��L�K��E�v�ߡ$�o���]�D�//
8Y�����w9q��N4"���~��� c\B�X�XƥF�ؕ����'�S�ݗ2�c��NBUnw��DI��Z&�x�����l=q��I��a�s��c����PK9���?T:�|kh��)�pN���k�E=[ɔ��*��	��,5w*2F�]1qj�f�1=#M�ˣ��z���o���e��?�^���^@K����H�פ��&~�O����j�P܈�b���G�����_錰�y��%G1U���k���¡e�p�0;v>~?�u2�#���y�Z&7�3TSGp�#�ɴ���:r!I�i�,�u-�f9�%jD�f����&5�Ickǔ�T��g�3i��f�$�8�Zs�L����"|��2��-���
,� A��@��Pn��w�}�b��� Ӥ�|(0����.;�f��+n���xO4/��m���p��(�v�%骕L����C���F{�	;Օq�u]@���<DB�b���"^�$����T���?���{JZ��"__�N�%��mc�׸�-2�}��T�%ϯ�A\$B��G�� �2�����|�l7����6��g5s�8MHE��Ziм������8��0�D� 2�J8ቬ�3�+�K�����*8f���ǆ�ќT��ٍ�����d
���k⠟��d�&	E���dcg��3{ʇ�{�OC��1�M�^3cS� E����0����xX�먀K�&;7�*+��Xv��+R-���%�_X�B��YB�n�us�������EK#|o�Z�����S2)��.s��8��iݶ
N�� �.�����}`�5o�
��5�4�P]b!�7�0�#���Z[ ��lT�v�d��o�3��)�]8��=�ss)yyZ�W���z���v� �mI%?Z��#�fb�6ܪ�o�d�L?�іPu0}��J���j��R�[I��s�yYO�r�?v� �U�e�����.�����ZIb�Qmh��h��M�ƙ���̚�'N�����?u��Y�,'JJ��;�����]��)�"k�����	�´�
}�GR\�`r��f{�4o�m�qh}O�7B��O��b\�HEyE5�!22�(�~��
��_K�b�q�?x@�)�c_j]l2���P;Y�?���H�9��>@�*5��1MȘ��~'�`�am�C�n
4�Z�pvz�qR|�=��X��#����U�����D?����&�.�~���7&�`ˌDl��i��zN�ٜ�%��%L�r���ԫ�� a�;#1Z)�mUDRe�Mh��c��f��e�R�iDP �
v�XW�����z�q�V-�RC�G����n���e1�qd�]t�����T����=RSВ��(�ՠ;c���a��ߤ�%�V�Ի�!�]�ʚ԰z�L�<�f��k�9�s5S��M@�? ^��)x�%ݓ�^�]Pn�p?b�ܽ���T�s��t��j5����v��8��rXE��N�X�8ű��G��ᗅ���闂�M撨��n罈�wq���{��WE,�q�z��0'�pI���b�����&����W<9���g�w"�k�.n�3�<O�^��ꪲ��~���4��r�%�8$�k���]
���z@�(?zB:�ͯo�܂�<䒁�<\ #I�y����叨�Ό�Ӏ�|�ߛ�p��4u���Kp�&�4�>s��yB(@nn�1b���&�h�b�8��4���ɼj�\:���4����!Dj�?��!=>��U�s\x�:߻���\�����7��y^v����\�)�WHԿQ����G3Ķk��RTA����C��k%Q/CJ�G�F�����j1^�b�`�kV�<V|�xu��*!�$D�~a�f���C;E��u���(!�D�<f�՛woߐ��*{�$�ꯎ.�yȨE������<�`-^�~o�l�
���{r��z��E�#&~��$��M�C�-$��	��y���i��ͺQֳCv���r��9^ܥ�*ժ!�TG:U϶~ł���!gp��]�ҹ��mݢ[<M�Ӳ�E���]ۛ�r�U�M[xQ����d�������3D��on\s�,s���aD�#�yj9��c���+|+�N��|Y��?V��1�-%Sr���W�.����o����#U+����r18�x�ߣڏ�<X<������">�,�a��\^��\���A����^m�EUk5�`����^����[�mIlHE/��Su�H���%���P��gtx{���Q�{��дX�E��)�R� ��䪤��n�"�S���ĀF��p�Z���y� �Kv��	lp�����$��ymz��+������S���!��S߁,l�)���=�㯨Q�Q|�G��5s��L�¿�to��uztjț���y��'sB.�& `3բ��b�����q�m=Y�2�n��O�Z5�n=���A�Y{8��X��E��#(�K�Z�6F�A*�8!�7瘢9�L4�fHv���̛���D�,��3��َd2��w�5��������5P.q#&.��N;>�U%���	^�xȨ�HWfY���D8������yH���e��\��hz�*_��(,K+�� �@�KG�Ҭ��s��O�/���&��*��m��o,��~L�qq��4��NA	v�ω��R��D�p���Z���)�� &]S;<S�7�ր��dS��F���}��q�~T��Q�VēV�:-�\s���3���Cݕ�Z���T�E���&s�#�N9А������N�t�q�e�����x�e���i��O��i}�򠞙�tc*�[�G����Y�ݱIP���j��?���;��Ӿ�D��ɛ���6͔z����i�(U��p^>�K�tq�D����FZ��pG�����b�Ky��>���Wg4��H�:O7H����U��j�t^�$���$Jg�"2�uFMuC��W����ͫwS�Q�w�&3���&.�Nf�)#T�P>��S�4�y?�Ɲ��8�&q�����&GN[��{;�A<g("P��Z�1�~�I��
h������L�L��E:��'��29����a��� �2T��|�����xy�}p�Ƣ�� ��7�r��o��x�\�����,���w@!�� ���p/�d֔ 0�l����t�@g���h���;���q�̸�N^�S>ęJđULn;T%������C��ߐ��_��<�!`��Z�j�;5
�l����hG��z�>]֕)�6�$����3��a4}�Vz��`���I���nӤ�G[L�x�}{a������3�@����O�m
�i��G��^ͼ�=0���XLU|3סtĴX�ք�_�xa��glz�i�x����J%��7U�3�v���\��ܸ��34�;D�{3�,���b�=0�;SA���KP���SgD��th�k�'�,#�ԻH�<�&��*�tz�_q���ɭ�:����(&A�x}3�r�o��.��!!D�/
f��0Lk;�Q>���e:�FAŸP̅�J�L�d#�i�P�E젖�؎ W�k����߹X��b�����п2�&�i~�sߺ�-;���q�@���.rG��T�<�b1 o�WA�!��z��Xۿ�8�CW�I@�e��O��Y������I[Rh�#�����^�;#�ҁ[TzB�>xnn�Q��-��u�p�I��;�]�������c�R�cb�=o,�Fп�����m�:��%��� Tq��۳2=eѽQ�g��rq�B�-%�qtODMUUΌ����˶x����d#�[��)h�7\�P�q1�G�V�4�s�^h!%��wt��D�����t��g�VPm�J9��h�Lp
�w��CdG,�Y��WW0�,�9��T_l�G�����Ǻ���C���y�L��O\�ԏ��8ĳ���*����1��f�ҩw8y|U��̻��z��ׅ��:��4�i�L�:1b*�����h��7�^�$�B�&���ӓ2k�O�S$T�{�*u�>�� +�P�M��A�!�=|wE,n)8�y��$�ܜz;� ��wB/3.�Ɂ�v�$/��z�g3'rհ�UQ<|/��֟|��fc����;7R9����ir4�5�ҌK���]z��5�c��}:��BP��"�/`��}�@���Ν(�cTS�����`���dֈ�`��!vu��P-z(]6��
u'�
8r�! �L�z�1��kg?�2/�2�2�<��I'��gF�al�wE@�y�ã��|vp�@�eBn�0R��9Nl��{��ܨ���ج�V~�X���hxx�n�:>���^�bK˂i����}�,M> hx�F:���X�g�g�6�Mɕ���^�|+7@�ĸK}j�_,��)�q*�{�sà}�>HQ��{��YزHu���#0�r�:�KV�KB�m�m~�nN���O
_ޥ�]f��:�V]-M���j�j����y*���j҃��hj��:�(8[Һ����:p�7K��I��=���Ӟ�Uv��]���0��3��4Gm�p�S��v�l ��#P�Q�A-6��VS�/�5�/yj.=�!nt����8�&���S&'��L<�B�V'^U|�C�Ye��(	QQ�y
��]=�e@���N�qSIڼg{d��Wa���p=Zx���0���<�������b���F��򠃠�^f)슈ko� �[>�����R����[�iWÐ/"@R��ۢɓ�6	C��[m�Omf�|��C����%&s�`Ґ=ₚM�;�Á��O�v����}�ǃ�+G1�%���'gn��{K��Y��0Ň��j)f� �^JȄ�J�=�m�
��EBI]m��)�f�R����Y*���u��~UC#��U���6�5d��Щ9}�&I��V��{xL�'����,l�����#�{�I`����`��%��KyC�-�8 ��>Y���(�C�t�;|�Q�]��L?:v�R������9aC���K锼IOU�
�a�O��[&�`�B�{j<���Z1�?��C���WlU�i��V�^-����-\����a�E��WYxZ�`2,ed���袳���.mG�͆÷�-�'XH�����?FH�6e>E�4֌�d�����3��MV,�R�޷8����.7����GdY�B�d�ؓ��{���z�#.?ѢSA/�Ӻ� �Ì��y����O��Q����P��rus�\�4 �9O�wR$�$	0��+~?� e|��ABB}>%Mgv
l��T�VE�&�c�=nt��~<Q�		~�֟�U�`fN*h�9ʘh1�XoZBnծ#�w-zH;+��B5.g3�G��	�}y�# ce��a��]zR���N��i��v"6_��|+�rL:��!!%����<���)��
��i�a��k�	"�j����«2�u�aD���B�밲�9m�P����p��1�Ъ�{:iK�:�z��柶��K��7��\�u&�]v����C�T�D����^�\�3W���}J��V�ƴ��-���>������hU����MZ3��|�۰�2��]X�ج�V�9��4H�B�ckV����������}!Ù=I}�����!1�_�&�G�:��-�R�8�,����h�� x�h�pʾ��ͬ�X�?�	m�B/\�s��^��+&�Ö�μ��>�Yp����e\[�U�n W��w�Y�j���C,��_����K��'��L��y����W#��}i���i@d��Xj��p�?ڕZ����:x�isʣ�%̦Ųцm�"�>�ZrzUOcҀ˒��&m�,Q�9��g*;�u{@�@����~��|W+�P� ��{�J5����3��>{�.n�4��į��#����3g�4<�{[?��4r�\��zRk��������#N�@�WYH�\i*�e�](!`���Hh�}?�70H?�o^�}|`�
x!�i��+{,Y�xÜ����S앦Q��K���EE<�©#�ANXW���'�r��BO_��y|��js�I����̈K�)3�����A5���q�;&�i�]z?��w�h��G�ۡhH�����Ⱥ��U��K1.%�S�*�CS�5�V�X%�\��i��n���4?𳜶��M �����·�/<��)n]�sJ�zo�#N1�톼�R�o��ǋ���T�E�28��5�y�to \��[ݲ�^�{��D$v�b��������L�0�5��!�;U9%r��~�zP֪�B�a�gu3�j`��@�u2�J�7�j��H�JVm&k�'K���E��HPj�(%��t�ˠ��2��$X��֓	�"`�9^�Ⳕ��U�e�4�Ĥ��	I�T`]�E�~��p�2m�&��^���J�K���q�(�����3w����lӭå4��]�_�ʻ�.0X,C���ܖ���G��-�oy�2b���_Ȫs؂[24O�: �����EB���iH���n�i���8xH�߃b�_��}�}ce�~`ݰ�$28Q��s� q�C�N��F� $�Iu� �Ƙ�}<��
���UmJs��I�H�~�t(a(r��-�3[ZO-� ��%8�)�����.?�P����C�i��M�ZG�rFL�}x�D��U�����v���)��}��%»uE�
�y�-�כ�$9�L/�P9�WB�44��8����r. XB(�bqIo_VՔr	�_����6�g�`�c �Ͻ �a90J��b�<zF��md˸�����!f�Yt'�l��;�Hٜ�r�R�KCs����E5b{1��9���|��h"�P���ʄ�{�6��z��nN@�e�أW�E����cH�]�S�V�(K5����ei��;�N�H��.�}"��k�������u�ɏ�+Lt��[��J����#��p�M�^	J����^k��ʵ����IP�>��;�Y��ȅ�3�0��7�����j�.L&n��:���8��˓�7͈г+���
h�����Ơ�>?�>��-b����1�<xR�x���rUt�xtL|_
�i�#�<ܫ~D����<��M&�HA���ԆDo�����2�
�7F�˛��	X��Uw>\8���v:�E�x!��Q�.Mi/�!N|��@��	b5�ǈ�}0}C�ɪ`�����MO��cq~;&�,���O5�Q��-��L��l���X�s����ш;L�9ww�:x{ �iRC��2�)�9q�����ңRL/w�'�^͖3��JK1��_������)ء����G���:�˻f �fi�_��_'9�P$`hN� t־��4���v�9�8j����$R�L�2�z��T[������>3D1����!Y!b�p���[�!�����t�e���^`���]��ԭ���(���T��tF�����yQB�G,²�!Tr@<b�hX�����sO4a�n����qI/�Z"(�%g�x,˺����n.ͮ�_�D�Č�b�tfq�\ Z<���,���3^���(`jN~��^ζ\T_r�ϳ#9�N>3���ӽ���a#4wrnH��˴۴50&��ʻ�S�� ��q�`�[M��~#�t��
�{%K���@��ɾf���s�ľ �Q�z��(fjB�~���B��uhC��d"!j�Z>T�n�X�5r�-���^�X��V��{�&$��>�c��n\���˕���;��lP����N�s���b�k����4��H��ݙ�%Tr����W�bz����m*�R~
����L`�L��!�ݔ�a��ZU��:Ӽ�5�L��c3$0�1!Cу��4H���������V	��Ɩ��&垁T��������Uw_ߪ��E5$��n̤�6b�>�sg�w���r�A/:׉S�To6U���F�`]b��ڻ"ª0�~����jbY�W"�g�B5&۔�My����MD��QM���������0�u�;3����������RC��4�&o�؁��-W�{o_J�Q���@Z�����{������-jSȑ� ~,��3��Ch�DT����{H�5�;w^YU����u�5���W�x��?�ǔ9@�^������HR!��\|IN��툾D)�X;��X�0�c�x��t�لڡ����L�[l����xr�cz�]`��>�$�oP/�޸��*ψ7-�5R�d )�_LU�����3R��1F�k{%�InSP@�F��I4/=��5��!��I@$!�zض߶�9��?
 ��M�)e��z�i�;����]�e�ޞ��H�U�[0`�l�����M�$R�$K���A3!�u�� E�Tk	GhGl�m�^;[��z�I�$�$�,���)���Q[5�^�<:%%!~�I2T�>�tX�Dr����"�4�k�`�7t�D�zmb��26h@�$���)��4���JȤ�ҽ��0� ��:��p�Lj��bڟ�=<Kױ�(z�@�ŽL�{�h�8X�+��ƚ=��������G�c��mE��zmV��r�IU4�\�
�R��>g�tp�MJ4>���k�;am�������WTg��<U}bD�vE�N��4ӈ�x�~�M���[�޴zW��>�7s��~���\�;LY���SLX$k��J���:��i�2j�5�����σ��lꖡar�@z�5 ����	\�#�W�/��G�5�!fˡ��Ǥ�2�I�-;��z	��9g�I�$le�K�t��h�����׺�{��NZ��Dw�mj-�$6͐�
�֏I	?l�����k�s��6gLb����#m��o��1�;�?NYR�m:�B��ز���ǐ��mZF<
��Ұ0��+�<������_�����_����U�y[�����&�$DaJڏߣ��.R�C#^����W���oi�
-ޙ� ���ǰ���y�
k�� Ȟq�j:s�/���/��<������j����+K�'���U�&�������wF+:�VI/�t��2����m��;D�\#�_p�>��v;"3nG��Z�ᛉe$����&��o �*Y���a�4�HנP�ԎP��ްl��⫡{�e�i^�(���z��ޜXI�݁y���k�HN��pD��r�e��;v��;ڢ(�
��� ���l��]�Uk�������ۢ��F�dJ¡�t��{�u;Ak���a�E:�z9Ƕ���2�ӏ�?.'��v#]�ã�d�����d��Eq�(ʳ�fء^%r�N��Y~��Y�>�&��^;\�7���h΍����茮�_�߻ٜ������~����^�D��2t�e"߆tuF�ޜ���Z(���p"��}�v 7Ot��H�7�Pϖ����Y����ż<k1�Y�R�߰}=|��X$Ô���b�o�8�x�Ai�Lr m������5�le���Ƀ������}��˥hW�s㷀nVJ)�㴉"(/p�����H�𯷱�pDyS��XJ(��c��OKC��9d������"ő���|N�����C�[�sz�Ո��j�m���5���2X[w4����u�U����k�N���%�MU�� |"#�?���B��F��J��~7��T��p���`*������o�@h)�QiѮ'�;�[L�B�-���\s{~Z��.�Q{���,o�l��gu�S�|X��\M� w�Z��b���?���=�pY]-OM�k�g~� �$��YJD��b�&ե�bI�B��A̬I�d�&(�jd����X�/߾My���.���B��B�t	e��e�9x9�c��|��I�P���mSy�i�i�V'r�?��7x�B"s�Uj:&�d"��NE+q�b�e���/��(%fb�<+L����[M����.вJ~�.��$*� ���^��*m�џ��}�p��Ȓ�c��s�{�P5�.�4PG�]��7J��a�/�+?&B�8��l*�����q���1}�{�?�u���d�Q}�����|3)��B��ת�1�]��?�­dAmG#;�gd�?ی ?;$y9.4������S��\I��5���H]QW�(�v�>��v=�2n��5�R~� k�c�1s;
�"�*q}�|����X����;�`����$�N�#�S�҇mz��-�>�ôQP��]��J�a�	u#�*5L"σg�Bxn�+))�-k���b�eXu#=�A"�w�t��q��H���FmR�v�z�[��=ճ-M�A�LUwY^����β���:�~����C��F�/�s<���!�3r��Km�p���Z�/M�*J�����0$�Ϭ$L���}�E*�(8�M�:#2�ψ�9G�}�C���.�+��!]���1�ͭ�W� ���t}���~���Fe2��l�;��r���_��p����*Խ8fQ�F+�J�=ߡ
��4��V�P��sE2[@2iĵۀ�pD�C�l�b��=Č�n�l5��ʦ��#���/+ڷ�iNR�D?�����&�`��9������uG2&�>1#�����B>�L3V�X�[��z����3{nD���T6���j��tӈ=�im���j�%	����W���A�
>�Mי%� 1)�]D}��OQn.��?����9k嚲��t�W�Yr�~'v�{�� ���bO�c�\��&a� ��7��H�r
��vpn�,�X��������`����H�~!����ydd@@Qk�G��~JF=�(c���,k��V
��OnT�*�0�z�eU���a��B��SIA�}���C���`����j\P�gԱ��5������r��R�{���s�ZL��e�^���u֮I$����Ely�����;0�m�k_ќ���*����HC�{k��n:N�M�Iuu��w`�xMd|;ه����!����:Ft���O�=`~���ɮ���7��(z�'�~�Yh�~<��p��<��	�v���q8M睌�Ը�N
N+��֋>IͰ����)%u������iAY�됱430�f��/8�+SFfI{�eKF8�<0��_#0}٘��*v���BVfV:I%��a�>�^&3�Qs�5� �:�����8Y�[5�_!V���S�[��<ϦJ��S$ǉ�����7qbݽ��O�Ȕ*�i�Jl�}'�	�kw(���H�&���p_< Ge�_�-��IJ*�Q<��ws����f}*�!��|��8l�f���9.��} h_j�Q��˴?SIoa��
]$>�Vq����6�x�GBTeA�:�w؎��ЍK��x:8Z_D����1�$����V6D��'fCLP�Y�߃��#I���� �zi�
d�,N^�����+6���:&Ю΅�6����bhۑ�}yb�J�(c�1������������耶U��_���4uB��1\U�m&V���:B�<���X[��>Քw�X��ޚIV��h�m��	h�n>j�+WJ�`�� ����'v�Y�b�&��������_�b#��ψ|�OerEA�#b�U~�O�L�,(���3��L������6���Q�X�^�S�+a����R�*si>N%9����*��m�+g���/ B��a�I��Гo�����VP�հ���1T\?�v���{�6���a��A�Ờ-�U�zO�(:��}\4좇2ȉ��ҵ�c4#�]�A��RT�u�9Y���E��u(�5�Tm^�ˤΌ�	�vc�3�h���T�z�y��u�0=?�w>����ZS���\,�2#�2{����&+���5� t���F�t�lC�XG��_O�U�G�×Ub�bVɀ��AXD�T�^x3d�D�U�jX ѝ���w�Tv��gY�F�MD4�v��
Ts���ے���d#�ȿ}���Tپ���KO;	G�D��ENv�>"���dԮv�j����+�[L��0i�	�a�G��Dߖ�p[ӿ����4�g��Z�|���IPri&�ľ� 8:���8z����KY�`'��}3F��6��ό�g0WpD���С�#1���'a�T-Sȡ��J��N�<aP��y"��n�1��tI�����!���b��t���o���C!g�Ti$��z?��A����`�u��EU�1l�+����y$m�i:��M�����/��I�<HM�jD�3�卐]�3�z�-�t���
f�1�z��eM:�$,��~��u̳�Y���ë��=��>�N�3���.�2��9R��zhnCl�z:���tIN�H��t�����?츩.f���?�:Z�����f��{t#�c@c�ɴql�W��v�+ �F�i(_����U�C81z�(�a$��f�H&��7�:����Q��:���?�Fr�U��d߸���1�}�C�����x��U��� �8�\n=}"����%:�
^F�q���`�qB.�L�䱔�F��Z\X8����NB�I��7��J�5o���>�Vv��r�cR��o6���H�Ȣ,��V��Q����	�G�,J���s�VI/SyΑ���"�D�9��S�0J�t�aL�W �����z�e;��.���7�<�$}l�1����X���Y�"���La�����8l�_�0n�b�C�߬�oC������'�����W�5[7�.��Ng����c�;�r]E���2O��L8�6�|�IGj��j�1{�~�Y��<r�:��d�KrGVA�|�9Ee���U2߲���y�Q�5x΋�i���u3���#�#)�QA��g�v��\.�K~`���\=B��7:
]C�k�Eq.}gH�b��\�
���%���]d�l������,$�F�-���׎׀缀��l�Z��F�^w��%�E�����4��(֡w�~k�{��U�O**��\v�ѩ2+#a[��D�������6�j"zl����S���}q�I�K:	��[���w��	�;c)��(=2�i9��y��.ߍPM=�j�\N�I��q���m��l�nl�"jjծ�)��� ��#��d����Ƌԕ��ݒը^�Z�-�I�c	A��;��4�m���hpGH`h"xiuQ뚫��a'Eֺ���W��ail�S'�{Ǘ��@Փ�<��P�,G�Y_M�e"�8�����|=����	a���M���],[�q�z�W7))R ��H��D�ɀN��y��"w����n��J�aJr��݁���M��9M^(��G��������f#�]M��;n=��'4/]_M��ғ�݁�g�fT��L/���]q�ݢ|�)��N��p��i�<�_�2�)Ө.6��,�Z��tc�k�W%
٦�j�7���O'*o����f���.�H�W������3BS�T��A��&��8ڥ�wP�K$�bS����='��~c�;� 0<��i_΢���^��].�/�0��D���ǔ���xL��!��$3{����,I���D���o���&بh�� 
�����4�s ~����z<c��	 ImH�[}E&)*�Y�$������_��BRI�Yںz̳�'t2	����Z��.�j�J�)h$����o�ވ���:8i;�m��Y.�+i�G��*��@������'����gX�޲�hob��Vr�y�����jy��֬��A�o|�C�Q���pL���%.+���wD甧/���#�_�h�Ja�:�}V��ꃧ`��ɸ?�kY���ިZ�b�Ӥ�m���,����b����YXnS��t�a�M��^9i�
^���M4��0Ӂt��$:p��|6p�c�#����f*�O����E�ۘG�	�H�,�AwȶY>�!{����Xۓk��8��.�a����\�i�ԞU�c��Kb��Lv�*�L��[h�o��ilLCL��&ra>�Qʆ�꟮����=֐�Ȍ��y醹�.��8�z�����ؚ�|�6*5�؅g���A�"=t�|���=Q��.B�d#.�����"�T�[�8��B�W�+���#��0j6𰎴��O(�S'?� �i�RQ,K!�0X�w��b��v�J)%U1ݏ��!Q�Ci�A��8IUجc�l���i�\-�l�����l�M��gM�$���k��E,J����2����DJ���0x�
ԏ��Mh��K�����'����p�b���`��\�h�+���8��tQ��I#�m�ބ\��UW8]�w^ 9��J����׍Y�1�%,�	4x�u�28faNA���A	���E0��K���h��]��p�d��,��o�2.�j��
M���9��E�N���
������4l�Ay=�z���DR9���� ���ؕ{���چ�Z� �:��%��6[�M����'�����l^>Cb�����>����{�]�̺��7^=�8!�6y���ih=�����j��2)'�x%P�@>!T�X�,�(-`qd�t�ïz�b5O�VV�9&�bs=cd1Mo'�	�%��z��:�0���c�{�#ɏ!�8�v�T7�+0|ʞ���K��Xyf�)�w�������0K����bX���Á�fa��z�dE%�1��U���
3��;*>A<q��g�A��H�P��e�����C2����6��$Q�@z� ��D8�fr�R�5��A}!:;��az����-["ĀG"��g���=:�IS������4Z�+c�sBX�aLK�)����zD�,�[�,Vj֓�'�����v��ܟ��2
�-��İ�苝�W�Jq`�Z�"����a1=�Kgy�
]X2vTz=P� |�9�k�~úm�by]���+c�9��d���^{:w�q��e���H}ΐ�z#SA��������#��Bd���ͺ����z��ÙU���N!/Tғ��Y�Z�~2����a�1P�"�����ե@h)�&򚺋 �L�p���/ƙN7̩�
z��U`���k�Q,Ȼ�U�*% ��xr<�[�X^H��L��ʞ�/˓���I���z}���� �"�'S���.Cg�go�������W���-ȉ?���K+e2�=��Eh'��A-/�%�;\�g����F�e��3Q^G�Q-uJs�u���!"�$�������φ��f8TQ][9R?���=�3i�6�K�ą����1�}�f��w���"95l�Y���2>#t�Xo�X�qa������>��I�uMO�@�h��9����/D��!c��Σ��-fljq٢~o]-d���a��*��8��6@���3�xu����.����F�y�u�H^M$�����5�!ȝ��-�ثit�E)��GP����ݾy����f��ο�R]������b���cE��4�U_����e��]]jEɍ�O�_�pwy"�,�~����n��?W����J�I�_p�e�+ L���i^�q8��iwO�Ur�[@ҵ�kh��8��)J�#�������G(���9D琉�^��L7����9�NoC�
]��w<gܴNR;+@��*���i��%0��⩲1�o��o��_�-�"���<i������h#��-(+a�������� -�9����^��|r5�h���YZ���m%���CjT>�/V G�>����~��c��)�Ӣ�Z�)��s�Z4�p��?.O��FW6v�:F�1Z��$��j����rr�rΛ�Р��B�����������qft�<g�Pou�m^_B���4��8�`���C���$=����u����'�Fш��-�l���:{�&�`�҆� ��f�k��Eu�|%��E�	�7���*yZm�eRI�"J�}/��al3�V��tp'�;�8��;Z��M���2�*�S��1� �b��!)r�z���a�j<ObHc��k��{sSf�t�a��j?�3��]|ǀ%�e�* ��c��A��CM���$�!�j-��_��m�;H-2���^�y܇�T.NF����j��c����s�t&��"��j=*�of9`���;�q���uH9(,�3�Ms����W8z����`����B)PB�Y���֟�&h��q9h<^�p��Ruz(�Ǳ�+	��:j�N^��T:��`Hh��j�f0*"1�e���d$>�~rk�}���l����}�"FWZ�ib���z�qM
+y�Sƀ�Rc4�'m17S���Y�wx��n������_}KA�ٷ�����-��>�W�T�"��^/����`�g�|@�N ��|K.��*��(W��K��Ε���vj���:��b"@�{��E�{�iU
}����l�K��K�*���$�Vޯ�ƶ�E۸�0h4����qw"=���u��UPS;Z�v���]d��u;��8�� ��Z� "t� $��	�M������>�~=��T߱��Xħ�'{#x��t�3Hv�n�9>�1:!2����D+\��5ef�����p�`����dNp}g�]�<G)P���? �SIT��ҝ�0�4ތ���Gr
y3.����$t�hMU��9o�[��&f��VDJIi^�>��+}�Sy�������m՜��h�d ������2]�:c9d�'�hUw焿9�Tj�{������B���MaG$�{�n�B��} 噤=��>�gU}A�@@���E�?R��3��A����ÂE��R�5͙�����ж	يtYz��P&�|��z�E�Ɏ�t�v��fz�h����#��/Q��k��o������L���F��ܿ�-�KD �p�-H�O#sp�lͪ��E�q�'�ѡe9��6�r��B�f��K��a��IL��o��n%?8π%ؑ��;k�&up����@�;�f���h�иK�>@�p��	�o6$2];��|�f�?�� ٱ'Oʿk锃���2o�";b0(�0P�����lpK���O��t%8SB�Fό�\���eq�z,�h�Aq��&�s?�E��<�Ӳ�j�˅lr��� 8x��G~�3cD�����4D�H��c�˩��VIϘNlM���<�}%L�������������)�)� �!�����>��I{�	�u'Il�5a�TC��yؑİ�ST��z�&f���"���𢪄{\����Xs(P�Ŷ(�%�"��&$���J�iħ�g��%Ď-�]���"��'-+��K�(�1�6��G��e�4��a�vXn�ͨ�w$��ΚrE��Z��f=f�T��݊�Y:�ZZkۨ��|%E;#��&���8V��7lz�\�h�E���w�U��`��OgJ����sm��Zu{�K�uy�XoO�6�g�_�|4ɩ`��V,����5�Z'���ł<؍�Q�k�еÇ<����(:��	�0������9b�/ ��E�՝vC�-зM�C>6s�Դ�$��<��1b?��6H�F��q�����@ jZ%�f�h"a�NYH�`��{����/	�qQ%�J�����iQ?��i������O$�m�4�x\��%w!/Y�3���^��c��I���4I�����.*�E;w���E�uck�8��6{y}�LX�g���]P���Z�j��ԦR�4�/<ɼ�q��`��J�Á�\l���-T	MVwî�{���,�����C��"� ��w��P�����ӹ�aQɖ�ԍ\\�Ip��
:`])7�$Iկy���f���g�Wcؿ��Y;�>:�}���q��/��h���|�;�\��3�!ɭ�FT��2<Z�Gb~�G2�S�]�
��(����7*�ϭ�V��j}$C��{F1�0A^WS��S�$4���Q'gJ��*��IS��cw/$�\���
�^�-{�Gj���0M����m�b#,