��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w���>��!S��'ho)�ˆ�v󃜎�u�G�E?! ^�ZY�����m���<˨[S���t�sp#�5	�(1���{���ݶb ���Z���������q������Eő�-U���V�||J���F�7 ���gD���ș��-'���r'�bژ���ƈ���6� �P�>�����󭝵����쎊*�U�#a�'����v��!�5ן�t/�y$����D��7ȥ-���I���<EVk�M�ְ<��R�f_
v���K#�� �vS�����_��p����~�8����Yؗ=������}��X*n�4ӎ���ғ^>S��zhc4�����H�%�Q>��N�~����j�_p�"�'Ҕj���2�	I;�
.䐳b�:c�u��X-����G�s��ZL1
�R�`��B�NL�J�㹸��s�;��6��ӡ����Zs���HX��6I�[��+XVS[`я�P���(6�&��J 8U�چ��e�8t�iI�u+\]�1q�nrj�iߕx��l����O��W�v�sT�z���Y,�n	Jh�ȖS� �����s>}>�󏢐I���	ihv�ܣ=5�ڤ*���P��mE=�iI^�T|��.��QQE�_�s	p/]�N���D�i[�C�����Yb���:R��[d���RW��͍TS�;:^�W��hz>�>x�[|���:+>0����u=dB.�b�H�4�i����4\�Ȣ� ����EH�f4�΢hoI���1���=9EB��)U�G���	����z���$�J;zC�vm~�����F���%	:Ma1_,�
ٱ��z]ZL}��X�X�! �F�C�M�?���	�,����H̽�;ȫ_�^�9R�z��R�j�&e�HP��V��J���Mj*hsQ�`�ǋ�}��nFhSQ`M!��л��HE��.�ط�N�fܽ`����Oj��9>IDȨC�
~]Ň��ʵJ�V1y�͞�M�_GUi����5���?��y|%#z�W��)�\�@����|`� "��`���u�X�/͜�W��j�.�g�iPD>FS�~.d@��D׌ �OB�{��m�O0�V"�������P��'�����eƾ�z�`��G�Hin>��^	n[C����xX�<6#��3�)���ߖ"%_�5إ�v�]4�4yѾ�m*J�����%��Β>���o�^����c24tE�^(��x%L�����`�<�g6�)���;��Պ$����в4(*eH�����Y�~�	�� �X�ɖG�^)8t�	ႄ��V�ZH�IH^�";AǛ�HFʟϥ��7nX�Wc��q����1J�G��z��R��O���u�1˅����F*!�c�	�?Ѻ%�5�Z�&}f�9҅��� �>Smb��JX	�)��=�=��!'ʩ݊�nNG	)ck�p�m���M��ܙ���G;�������/�q������\K�o�jO-�ب��es(����~�|cC��/�0�������ҹך���ণ\\C�HL�{���X�Ic�${J�|��a�N��� n�¯;��.|P>�ٗ��ǤcE�,�k�8;ln��j@����#��l�A_d����	Eu+$�M�z��dk����ϦPW�<\
��&v�6[�
�C����,+��0�O�6m���?���LԵ�=���PE}G��=�X�ѽ�}��}J���l�ɝx�3�gB��k��E��3�P������n�զ`gwZ�-E���)~;��-�j!�;pyt�����J��Fm�lE��c=`���ۙ3�q^�>Mw%b�_��5X�0�V�j^�9���BA����>�o�w�չ��NP�6�0�.x̞K���	�3��0Y���{X`��0��٬>b�t�6����ܜ%e,��/
eá���w��<N4P�&�-�c���8m䙺.�32z뤘�|�{�,T���X����!D�ٙ�f-$h��Z�0'����/t)�`"�j�V��~/�����&Dقa��i� c���{>��1T�+����8�d�o��7�"~Y����sN��)F;�ŘIW�F���s�3;��<]:PZ�0��B����|�[O���yY�e���g�n�cj�	�E,bccpn)�Z� ����� 6g��||0���Y��%W��QUYq{RUH�j��K�PN�f*���|�"U��7�ю�%�<)ȯSZ��"~<{����L�Z9�0�� ���j}_�FI��	z����=��Q�$"��{�c_nP��Cl@2Lf�����m~�-Ӵ<?����3���/���g���G��"��@퓛~r#�����Bb����n��2x��������'����|r�q9/�����"�Q�b	m����)P>���\���&�s��~flh,$�U5��iY�~1�u�|�|��`�{�� i=
d�h@1;c������F���̾���ԷE�p�G8��.�;�`c{�����Z�朒7*彄�k4�ݵ.�Z-3����Ъ�`(/fc�J�J������Ə�3Ѽ$�%�-���d�ȴB�Ik�)mb�Bh������S���n���ښ�r�]���e�).An���u�
"aÄo��nQ;y�QH��҅\������������b�I�"WL��^�Bi�糭5T�O�︳?�⿸G͚K��hx�<6�A(���l��$��Re��R7�i+uX����B�w�s��<G8���u���+�M�h�x�O��y�wj��am��n�M����'���s�<qBo��$�5s���S�����KNi�U������p��f%~�Y��Rp� ic��i�����sJсw� !S�o�D���v\G1{z��/t�tN��;�%L�������Hk�V�$W֟���	�cT� ���?������$8��"����������b����-��G���5�h�3��͔����ϴ*�L�qjb�eV��a�q�����5��gecG\Z��`�K*q�����V��B�qe$�P�0���F��,Tqt�7�2�ZL ��] 3Ou��t��Pꕥ��/t���l°~fs(!�+�[�>�������[����C�uW�����ա�+��-��7@�RsS"�eည��|o�C<�.X�F����2 ��.
��_1���{5��r�lJ�2�c���?S}����Cm��s-�9o��E4�������*aa��?;زc���+P�8*EA���4�qV-.�3�H�i�c�� ,SEQ5���QM��n�g��)�������^�Y�Gۣξ$:�T��� �� �Hx����vi�v�-#p)��ԣ���}_Ŗ���I�t�S�I���o����U8���sYǸk�lLͱ�V4���/nZ�u��U�0���_��DVQx�h>�	Eh�]���ể�MdNK8����ָ���hC��υ*}��~> 
[u�� �;qGTI���-���h��{��Gߴ����S�ͺ���`�n��\(x��.���FV�0��7�#_m��f?�g��G� ��3tv81+�7!�y��Vk� ���e1\G��
[g� ��{*�l��H�q%,{ʙ� �\V@`�Z����'X4{s�J�Ql��}����P�5|�Z��_�A/�����D���J��Va�=��hI�U;�'���px%�� \Ny���bz�*�