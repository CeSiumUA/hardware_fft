��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c� 9o��|�~�+h�PjA`�z��#1LH�s6�"���Un'��jg�'g��xwaķ�E�ҩ��:�:K��� $�;a���9�IOVy�x~Q�XJ-5<^Zq�gr����l��"Y=%�_�����`%��t�L�"���`V�\�W٦�0[�}t�T<~��3�;��esJ!���/�N>=F-9���/�������a��H<+�!�P��4�懊���f��ܝ0�B��Έ�e�\�Sw�T>FB�SAن"`Q�IJ�~�ث�$>�]|(���+j]L���C~g9��
��
")��ֳ�|$�-SҨ�ʛ|}`���x
��ݧL;�a`�5�ܻ�������� �U^����<�����Q�Jz�.��엤�d=�t1S�2�fԚ��44���N�۬*�A"^|������7C�Ս��q��@By�~�ӌ�����~(FF a�N��-�?X���XqI�b���X�����l���50�U���!Je[F+���������4	~������F�����4�R>)�h��S��l�^��Ɔ�E��+��B� ܸɘ۶�S5����Q%�P�-��;��"��K���zc��&Kl&[vO�$F�퀓[���`�c������K1��q����O*�-�iN7����ޏ����eu�!R}F��i��]"�er�T��X����@9,Ȫfώ�;�A�>��6�"}�*�y�P����E2O�7�4���2�!�^����~b~�]�k`�1u*��v�7_��U�9���Y����=�x>�~}&��D����d����	x�����l��艁:��ZEGe��`��YWu��]1��a�E������nU:��]��yL�l��UN�f��RO����٫������i'��I��/�%��ם�k��u��r�Z����Nv]�S/��뫱u5����l3Π�Ӵ�$���]�g�[9�KS'�
�?t��=hX�5����_����[W�9��N�G�}�����E1��	������Ԯ��6ˮ�-�0�?L)Qx�}8�&�~��ݖ�^�6�����]�jG�����ʒg�^�W��:{21�� '�8�W��ks���� H��Vlp�\����Zu��'9&����糊>Y�z@3r#�N��kn>3��U�y�oq"V�֤o��]ۮ4p<Y���'��A��������F���< ���0t]��0˱G��7�Y\�:U���h�/�2���j&sV,�?�	4����Ƨ��"��	��$9��H��+ׄ؊줂_��b��v)2� �T'����^�-�|$�7�6,s$�l���UGl�l��Jo��er;�����H�[�tϠ�8F�����s�#�fȇ��+�P5���2���q�]�p�b����U��F�9��mr��|R2aW���k����t9PA��$�(`�����'XmI��<b���pTB����)�7zs�� f�sb*����[��{�hKE�����Fu�>l��~��V������J5GWi{!(S��@�J'؅�FX�0�Əff��=?��9�ρoXL7c��Y��x�t�|� �`Az%o����/�c��	X�f����ܗ��#��W;@>G#���=H�1tZ���r'�P�cw�o��-���XyĆ!oZn ���0I[Aߒ��דR�rL<ə�`�03���פH�HW�֕I���*��������t�4��V$�C2n~�-����r�9�І]���V�pc�.�S0��2�YD"�k��<�IG�\t����sa��33�!���MGQЙ�N�#A��{�k���	������}�&�^褿a>uE�}�!�S�C��F�QN�ݾ� "�N��� !\�!onl�����N��i;����B�5�,��(1ˠ��n��aެ�5��fL�J\1��?�p?z�� ���fM����:L�Xr	[G�~(�@qN!u�*�<?��������GV�>�=�]���tHݾT�"��@�)���2�u�K�؄�N�4.9��!��/1������1fc��jA��y�+�����~1��}4>-Md6V�CAv��"�K�,���K��Y���G+���?���� JTx
\�e�K���!��5
tg��-z��u:#�w�J��]�rc�Ѷ2����q�5�)]Қ��|/}�����յ��ă:��O����P�%+�HN������ƭb=��k�_�K�N����]��w����*ؗvi\%��$G��L��#H[��$�`C�����`=H�Ss6R�QY�b-'�����s#��{�h�:e�vl{kZ�e���, �k�e�
/ղ����@��@o��e-�R �2���#:�ÐY�����!�H�^FI,���`��4[��.4 �B��1 ��Bm��A��
쭌z8�R��c��y�Qjj#�G�W/�VB��=WV�]�9��d�V�$�)ڨ�F�-@v�4+K& �V*��I.0� ���g{@c�7�v�������kꕦQ����\��愓����;����8�^�\8��}4v=�#Z3�[&�i�G~ǸV0���T�L��l��3��g�A��-�gW6w�MH���͗v��q����T��)w]���rL �N'Һ��7��,N
�E��|eekOgK\�]i�]q<��ڔZ�E'is�eh��p��^/Wn���%�8��C2�oWѐ���y���c��]2g燺D��Z>�'�(�0�ƨ����|6I�s-�3�
~P�%�&!
+Nc�~l.���}!� (2��	�3��| M5��y/7|�`�R�_v%#����T	-�v�1���K|��`�/V�:\Ǒ���Py�J�VC�oǵs��a0�B�Nc���$��?S���O$����GҾZ7���ey7��ngNļ���cn�E� �6��ՃE��-���\2� q��XϛNS��z��q�(Q0��@	�^���W��D5�RM����آ"NP���(��{FS+r%}�[�����'�q���^1�D0��w���М���p��5�5��t���z�l��pQG�6~�Z��j�j�8��3����V�_�og+�2#�����3~�O�㒁���AĆ��U��B�����S��������6bT�Q�*�@h�������߀*S/��w�m2}<�>�tq��~�V�t��T:��[�\kn-в!V�2?N���hzX���7��,7���a�?���}�t�\�����5�L�a����;�*;��$��>>�(��Y�l[�g��d��w��t&���N-~:�-)åge����c�����{*��� Jzi\@ ��������g]	u�T�[�3:�D�̚k�+��0�+����U'�-��u8��'�� � 6�WpSK4ʗ��,O� ��&_��<�l$2��~�'k�}sp�3��t���U*u���v�V��.
\�Y�7a����z�-$��Dl�1I�H'�}�����~#30Xc�E�W����9'ԬXO���n�pG�g�9�Q1�9�/��q�\y�E�y��0;��R�U���1����Qe�fܖ�i���I�z<(5��ݡQ���V�I��<�6'UVb���C省 ;i���Hს�T�d{8��W*�8�s����ru<�Np�:�h]a�̈�^�&`���l��|l&��aM[4�R�J������:�bxq�)Ŀ%A��a�n��+Ӄ�ڲN"E�v����|��z�W&}y!⓯�wv��*2D�ǰ4i�p���+VZ���?��du���(�K65��5�q���C$���|�c�o:��miҲ�W����ER4��� ���17;�6aB�c�/`r=��F��x%��#=�N��}�Tw-�"��}���8�؊s��vRz��ys�Bq9�HD�j�SL8�X���K���'��l�N͕��	ڇp��P����x�j�`��O)S����W"����0+17�9�������Q�jߵ{Z�^�o�dܾY"�N��f��|3��O���Gd����GLnN1��]�h�oI�6�4�P�	� `,h%�ɖ�.~2�K�tKw���4���Vp�Cr���@s�nƘ���AKTD"��m�9�G�g�.)�U�n���p�5�u��IS���!�C���ض����Ɩ@*BK(����g �a2>I��b���l�Zk&Rfv�O����o�u�1�عV�d�#���޾�Q���1���,C�HS�7�E����l6�J��0��LNi\{�@E�Ns����.�^/��(=�i�׵%/xY��J���N?�j�ᤡmu#-B�$�E�x�رԓ>���+�3����7��s�U�]�uk${B*
ظiʼ�o��svI�7E�Ӛ�[(��oI�-�xby@+h���N�2�f�_3�� �g;����~�B�"��Z��A��RG�v(ٱ%
aBA�]��;wD�a�X	?Ln�4B&W�R��/R�boM�Ǜ��E�+ F������ib�D�Ӧg~�����I��u����T9LR��3��Oz�a�
����i���;⷟~F4�#��s���X�f��a;P��Vt�B_��Ya���z�!ik ����x�2�u�c�"�e|ԫ���䪤v���1��Z�'�F�WSQ�����"��Y�I���Ii�bNH��b�8�\|���~RП&E�P�z��ˇ�0f�S�E�"�*���N�V*X��Y닩���U���j&�_D���Be���U��%u�ʏ�ܧD�ݑJë��)k-�����ˡ����I �0�q��6���}�W��؞�G�!�{� 0˗�Q�IG&\�>՝�t�1K�	rx�KG�ڽ����.P lh�R��b�?�d �[��Q;�c��@�^J�\7�FB(/j�@Y�ׂb6� �	�^�sZ�L�v�T�c&�y���M�"�2�}Г�����2�L��[rMS���7~���:Z�"���Q��}6�L��4B �X����Z�ۺw{օfLva���<�?�P�xHF�$�`�e�]�!���{�A.�<��y�V���
�!������嵑���E���������W08G^i쥌q�� �Z�2_cb)��6%���pX8f���&�4��D�{�e�;���CU�<�%[Q�j1��;�"�D>[���f�Ѩ'�G[�,^�- i���~L����Y���G�5�]uO�Ġ`�[�����R�Rv�5��M��T�eT!bɽ�R�����ҵ�-�#~_/%�:j���mo�����˓�O�����Х����L,$��b��|a�N+/$��g��7�1�uk�B���fU�f���&��9�;	J5�K�}��)SbLp�y����\������3��m��vⓕ�ZY>�ɸ�����A���8u�����Ro6g?ibċIIyo1�=_�Z2����u�.B�s1�@q���j� A�k� X\k=�"[\��)��p���ŵY$���nN'�~If��ַRB�k��O��z��C��HA��rRt��̮�.x�n�_؇��l.��+�J�gJN:h��v$j5Φqli��c��#���x�� J<s�*	��&��J��K;�f��)+ۀ��y	�
=�J���^���[[:nǢ�<�� ч��iWOUr8��i#�-#�݆�A\3�	��r��K� ����eF�{OV��P�}�4���`�C�-��iH����iJ�ä�����]m�2(�
 3��v-�	�(���5eX1�6{�r0N%���]��a(%�>�|�Y��:�&�ї-��t���BJ�/�F�Km�,���7㖴�q����^
.�42BQj�9������F"����^�2t�ZV6�7���^`��0�*=F��<��(谖L�_ē���ڦZ�W�bw"�2�"^�w�Ʋ�.��[�2�O�É�?��l��W=Ba
�,������H���	�����еA�Blυ�/$;�SM�DH3�Z=�D���NM����م�Ij��}��_G���7� |�MDX|�gG`*L��%9�i�D�<R�9��Q������l�]�4	9S�7qU��2kX�N���\nA�S�+�-� A�fPg� �1�uˮ��JR�S�jgVю0>�9!g��
H-R-�O�352zH�_
�c�r8/4�z+�G㱜�St��;���Ia@�5���t\u7�L�<{�����d�yn*�v|.�f[fP|4/�����I��{�I��۹H�Q��r����|���-�	$ ����KY1���X��toǨ��ۦ$��~� �yr� �^�"t�Fb���>����~��-��Tb ��63���]�nA���d�&�!E�Eg��R�0!�i.�~k�kk7mU[�<�z���PW�ߡ(�-}@�Xu +Z:U{t𹶍��n�ɽH��*���J��� U�T����)�?pp?ݠȹrwjQ;G�*��~�Kʧd��$�!��}�;SL�z�_�+���o|�"�ܫF�t�q��#�D.g�Q�I�����崅�
.��dH_b&h�B>s�J�av�%V����RK/�`z�`�,tp���[G�}s!�R�(l`P�_�'�;:��	7g�e���������glK�`1�B�
�7��������櫀e��%�<�he���rza�#�o��p��F�P8	��¿[{�!)Xw"�Nu`��9��>F~���#����y�e?༦_�n�!٦�b�8�ۂ"u2���:�d�e%ib}�;P�O�{_�� A\�[�aSC�L!bo#V{1p�a�����lbc�35�s?�޽:��	η��s��@���c ��C�
g�_0幁F���.ʾg�E���60a�����o0�n��@p9�ש��Xa�E����V��a�j�Z�@�МN��l�~�Y����q�����Z\��L1F=*3H%�L̒>���h�4@��F�&�z�^�W���`x�����Nx�Jӕ��r�8L�s�x�%��v��՟��ݝq0eS?b� ���k� F�9_^�8ԃ��������EVɭ�g���Rz��ދ�Y=�b��j�aY�: �]�j7�,�����2N�o�vI�M01c��R燰*2խ�2ŀCؐ�F�H�]-�eB�I���)W�3P	Z�Ro�P�M����fǀƼQ�ZR,�o����J���ܼ���~��晗 ��o_�F7iA�.��:s��]�!W�E�^���3ĉN��C��i4F�;����c�#�G�X`���VBʉ�s�N��u�Ax�rO[��ȫ�xk�8鋜 ���[�rmSl=��Z�2/Te�֣'�����Mh����K��C�a�e��e0�H;�@�3_ڸ��6Sh~�A��OAl���E+�����R�nTzN��YQh������k���{� ^�KHyF��ӹS��]���⬤���;?u���~m�+'y�-,�ne1MV������3����G��i�s�1+?A�@�X�-�0����o5��ynz��݇C����x؜'S9A�M�6�g�2�O,aX�nb��P����l�w\�K�k�c:�[_P��z�X�1J�j�����h !��9�|Hݠ�M}������JS}Q�aPFu-�ub&�nc�Pm�W�Ѐ�k��t�:�._9�w����P��zθ���\Ե��B��c="�蔝��cݴ�s�F]@� �,g�t|'7�Z��1d.��dY�r�A6��/6H2X�P_�^l
Q��j�F���R�s�5��h�hubr�4i��L���I�S��W<!�12?��0P0���&943��]�d�X����{���x7���5�:�İo��^"I��A�̘L]o���M��h!�0��b�rvk4bi���ӌ�:
�	�,���V�7'�M����i��\b��{X�n���� mu��
���Qޯ���("���28��<@Qzb3��� ������������5�:������ChN�	��$:�Ո�a��+Vµ6*���Ȫ�\:��Fz��}m���6k��9���-Sr,�[�i4ICv�riB|\����i�`���=�_""o=v����!��q�>	?���z��\b�L�ߚ�8��ph�39,r!`�Ba�}dW�n����}{h�1FA{��D�}@ҞD�1��J��2��»L�m�	A�*��"����~�ϒ6k�7�_�+�?:MD��8J�~Q��7TV��rUޭP�$�}�.v�&:�)Tg����'~����a�Kn$*��sm�*���%'��ɠ�׉�$jc��N3*G��@&��d����e�`ED�����;�ݷP̰=�����jQ��~3x�Qr@/z��5�iG5���i�8C-�3�a�TֶO�_Y;;X��-@����F�50�( Lbv���P�ߑLv��-(��"w�]�~Zh"?F�j����O�1@!�<�;ώ���ꌋyv�o�q�f��~���1Q_hl:�L#l��1��jl�mF�PmO)���%A��O�!�&��m\B굋;��X�n1��f���Nz�"cc�V����^3�`�e#�
�裀������%;+�.= ���2j����V���MԊ���y~��������ƙ�
���ފ��{��p.�����G�v�8����:��E����r����h#$�3?��;V=Mb9��9�1��<�)�Z^���6$R���s6����CO\&}�AreɻL�or�3mƻ��ހu.�u)��;���$���a!"w��#i�<Z_�,rw��X������<�ε����t���&S�$���Fg?;ڬ�����Yr�xݘ�K�yv�ih]�8�4g��kr_����D�GJJ ����6fi��Uu�Cc��M�-^/�23^����g�1�N"FU.җ�2I,�A�;lhT��0Z@D�O�$�F���;y(T���]� ��b�8_k�7�:�p�&�x'.���$��~�}r���wC�%f_���ź�������3��Ρ:ă�)?�fi4w��ks�:jjlq�cױ�)!H�~6�#Xm3)�-��m�<��=�������ikp��%ͨ�J���ɃFʻ���ML���*��t4�B�Ӊ�7�7���F�Оvy~��,�i^Li���/{��9�,y��:]CH�a<���D���x��øD��U�]�2d� �\�h�m9 ,;��"L�p.�<9�b��9�'G�����Ӵ�pÚ��rJ�#F��=V/E=T��̀�u;���܁�S:�� �>gL�F��̙��П�"���aY�I�K#0O\N-�>�0�D�U���L��T�����宀[$��M��L]pՎ�����U���i�,u�j>�z��6�wvw`�T
�f�ńk69�]BX��hyI� ����d��XE)����޸��Cbٔ�~q�}6��2s�b)=3-��E��� �5�uk��6�=�������ly�1��Z4��w���n��Q0ã��I6���S�2/p�4G7�X�;P����&���	aE#z�U6��^$�&dT�8{9�r�a����'T�yr��B�+v�S9�
Z�aE�j?�v _�>�����<��d��Ȏ}�B�#:�7������vȠ���;��5M��F�¡/�Nh�	�Ԋ�fM�����meEP���T��ȁy��ܾ�;l>��>T=1�U�kJZ�>�E��6WRX5/c$p@��M������i��,����8��<�x����Č-��hU�/*�[��g3d9�������Ж�}��@�n�t�ы���1�����P?��M�����o��.IW�(���t0�� r�i^\�E��<>�w��<_@��x�`-�N��j�NU�%���ZޤYFk��@��qm��v�G�!F1��l�Z�1�&с�������%N�NޝF����f^�DZx�B�+���DA���XD�b��قO��,���v�<]�ێ�.���=ƺ^m?�
&NRM�@�{v-a�j���[L��T�׏�=o�w��(����Y�ܧ��KS�8���G璗���� H�k�D�J�+�e�0TB�U���=)g������p�T�F�@4�a�(�A�����ϘC�9�2v�Zt%
�&A�@����&a�:��:�%9����ǕE���e@r���f���c}���%����6v�F�f���JA1t�.G���b����]+��ڹ}$�>W���Y=��.>���]�W���P�"�	4�e>�)R��Ǔ�y/���$���r"*.F��E�S��/�3�9����i��.��̸�*�E�Ɵ�)�;:�9� �U�