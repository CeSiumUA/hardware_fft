��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c����������E��hA<�}/B�2�4|p(��oy�=��[�}+T�:"P�J�A:<N�gIE���@G�qt�?���o��]n�=��.J	y-�]���F`����?"��;�q'�VST����C����V	�����]��P3p���]��BlᏻQ�)���6��}��R�Jr�L��S�_D�-�Ͻ��T��q�B�c�$�b�	`jn>T�x�g[�����ګ
�Ne'��>ʭ�8G�$�����p&��dv^����8-7Z�|R�}[5:R�XpIF0M�Y{i��79N��G�7�j�$�j����oB푐ڻ�"�qPlR~�0��Se�-���e3g�e"VX˺�����L�o�w#�,!~Y�iG����@9�zJ�7Mo��.�Y�[�V�L��L���A���^�0���K�N��4Z1�3��M[�=�ܮV�;%��<9��'Y��eK��{1�B(7�RV�el5�ٔ��6����GG�)�6�q�4�o>+y��hD���i��D�����c ?3oI�+���~�7oi��ݣ��*lnK��S���e� �ԉ�7�/#K�FӟE+Ɉ�F.:ǘ�bq����_3�E�:�}�B?9@�˳�.~х:� ���~_.$��zhlč���ڥa�,@��	=h�k����NXes��㌃���e|���<4��0e�$����]��g����mژ��SݬЛ��4ts�Z{t��ŷ�G��#����'����Y�G#5Lʏ��0�ɝOX���i��˞��b�2�;�ML�r��ɴںY\����x�0��R�9yk�A_nX��τļ���Q�L	�1�DP���u�3�F�3�ŕUu��kׇ��R��1�*��a��I3�
UF#��i��Ł��.7��)Q���6B8b`n��x��L���<$�1L���$��[P�[��F�a�0+/&��m�6B���è�m�t�o���lm�(��Z��Z�`�_�1*I��v����9����N�� Vx;O������;�'~v�!��ţ�;�_��t�Z�L�M3�R����ZP����|Jl��0R� �@��Ab�$��A��Эơ�ho�Yj��ԍcM;�X������`�G�G"��������u1��]Y"|�0VU&04�j���P��d���(3W���a�����d�;bf�"ޯ��ݵ)�E���d� ��|8��KC��A��:��L��$i��]�f�:^f���?�WL��ǂR��!{b��,�,.p�/0Tg������W�s ,�o���ث�W��*Ǣn��n���1�#'s?\f��K+�*j_���V�B#�]_�c1G��ֽ5�c#�g��t� ��d�f�꿆��p̒����>��������!��}�}��6NK�{=��c [�<آ�2�ig��U1�_&�>V���Ȋz���܎�M�R}�EW;�	���m4�/�kx֠��]iPt�*	�<ػ�����8�n!~��y�cP�h��sr���G��c	 �NS��A%q��F��/gAYv-�?�)��`da��a���݋X��tR�Y15��3aH��յkm��RLIQ]��ZI�c��	mq뤮
B���R�a l�f�q��	
Q1�ڃ$�*��V����:V�(��沀�O���Y
4B�Klc�~�G�� ��ޫ��Ja���	i3*�>��i�JVbCW/ Sy9<k\f��	���R�:�ak(�K�n�$*w�Ks���LrA��Qk�������@y=SHQ����
��c�hVG�V�,FK�GtJ?� �Ғj[����T#ܷb6�Q<F������Ԩ�).=I	��Z���v�)���H�+a͇ȁ��0���7���o:��ܼ6�q�E(�i�]'�������8��l?NZ@΁��I�h��y@����4ü�����!F�����.E쾱�5P���eE3g`F�4+E�硌�$���	</`Bh���yc����f:��G��� �;���!��(\%5:��y	���D�W�Q�5��#�tN�m��Zg��d!�\8XY=c�.Cr�-�Nt*�'M�L.�q�}��z �M�z|���j<j�������D]�K�� �3�F&�i�eT-�4�z����Q�x|� ;�nF%�	�_��7��Ix��2=-�!W{_�>*�,[R|u�j7a\�|�G{������:*�|fx�:R�mx�le�4����X`�)�����!���0���6@eP֐�ι0��t#\����r �ë�9�h@IJly��Ծg����r�0ޱ9�a��4lw�h��rJ�?܄���3	��'$�fOgJ���O-R�D�(,,j��]̈z��<�X2H�իr���М6���a�x3��}��4%��WgX����U�ݷ�V�_yAM�m6��:Fi����.FB& �O3���Ԍ<WT%��(�<ps��0-^}�\!|�&�ʆ�^綞��A�Z�����\�+��������R]��J��wE
���'�栵nI��1���+<q��&�G���p{%��r���qu��p�l�;�`_3
�����'�ѩ�R]Y�ͅ�M��g_��Sl$�Ox&�������;�P*5��3�WƓ�"ʰ�l8�(ܞ������f��O���]ſ;�J�1z��S�_������r�q����W�}{�y�a���U�������L6��Q*Z"�T[!S]{z�T�*(�0^�Z�R�ޝ���G���^J�.�U��ˡ�W�@�'(�L=׼��7-�ʜ?av���\}A�8��抌�F1�ǘZ
7�T�?��{fRͳp�4јY���|u궕J5�1u�Ax .��T�M��M��L,Έ�hY���* �s��J���6�+����2�O/���쉳{ֱA�#١�}��H}�3��)����}o$�#�������^�1���ki2Lx?��D��(��eΊ+��w��I�G���u�5c��F4"ŽD%<��z`���>7;���!qf�&i�����h�o6ژ��v�"�ڵӅJ�8��ՓvztQDYN�F-��K�k)��;l^+Z	�P���r�*�r��U��@߄~T�)��Af���,��!��l���tZe�c���n��]"���Kd��<��Q(UAW6�p��VP��#S��!/����3!&�� ѣ�R_%_�?���ٿ�|+��=N%�k}<ZV����EqV([+�]z}~���U<POX����+PQ<m��s� ��Q�ًO1|G���Z���FQ,ּ/��Pإ�˓]Y��y�	�k˯;o.E�6�G�Nh��d��"#?��Ԍ�Ml@,)�P�23U��X���&{�AP"THmj$�K��Q�Z/nfs��+��x�XB�5���z�K�Ǹ�=J�'"�6�PS�I���B����
柼W���L�(�B�(�&�tC >�ӎG)�w&�q�:��7_�*���=���E���!)"x����.[�ѱ�b#j��\gKAǴ�Q�	4}�M�<I�� �Y3rN��YQ���OHM����3F���G�m���0�˔������^���y�T���[����&�'e��=�;�������qI��H���KJ���<�o�3K�D;�䥪]��/o����c�r1�;6,�+7Bۤ���W�J�Tg��h�bI0T45��{��^G=�\��'>��ji�Ax��5�M��=�m�<(/`Ý��	�
����f$�	՛�
mޟ��͜�̝ѧ�������17��E1O�M�澣X8����q��;�+��ȇ�YB�h�1leQ�蘛��=���L��t�un�QP �[-��=����*�����_�8�Q�/a�ߐ8��}[�Ϧ<���6��~&�K���%�|Ws��`�`�R$m8��Й=�ݡ��Tk�,$z�z��O]�/|h�Q���ɐ�覯3��^b�����e2ٮj`�8w'�����g�y�	nq�Uet��xǥv@�:�c 	����%D�o�ҭ�>�V�M�"L����n��Pur�(�g�x�ԋ�Ֆ�=���"ٷ�E �����h$ɔ3Л.�7%ɻ@�� <Yd�]�2S��gѝ�.I)ҩ1՗`^V0�E�`f��Ot����T�G��4�Ktx�i!���l��Rl��oTmY܉��������ɫ/��H>Zl���I�4΀�;�g���Ԩ`���xf�'	���֫�r�Զ�����&�UUZ+i�o�=��Jfs
�
��#zu#���<��f�]Ⱦ��<z��[�]��ܴt_�eg���`{���h�H˚�(�#�i�z�I��/��@�9�E��Aݔ�a~[JS;�h�����{���v�@���XvU�s����q<#��9o�����⪹Ħ�����<�\����쿰YEw��V�j۽��7��0�&��Vt1�D�Wn�ok��З�-��?��-������ �_��Yx��,*	?xx���S%g��
�뤀�} #$�}>��g�D��mB���0�=����Q�Q�M���Ld!�1iT�u��r$�Ŋ�ԑ��T��]5�+:G8p��4���5��چ�ǿ3���pp0賲�4�(�p��)O|˧��"��L]�������J� T�
�;��E�^�*�"�pؿ �KH ���������[�hY^C�܊��ߊ�eQNӘ��J��}H�����>	8�ҷyw�"�SS娛�*\���il��aU؎]E�:X��[�hS���=/�,�1M^�yi�N����z8�,�J?��16u�M�k�%��B�8�{@Y=�W�a�V*��W��o���aݙN�f����D��0ZC�����ѡ�Tϼ�:����rm��K&��+w|M����-g9�����Ng�����[��< ���0���y�|���hViv��yA�9Za��!@��_U��:�)�#�$�_��F�����5�s���������ۭn'),P��.����P1앗?�yQMW �{��9�Y��˞�9�%^��E�ȅۑ�G+�v�Hɪb�����Pm�zv�6"x��e�a��/�J�RdG��נJE�K�A��m����_P��Sf��YP�sq��N�S���59�an8!�#����t�^��v��f���B��aǥ���S��� �4��#	ۑNUȞ�B�Q4���[�H�Ԟ���QId� ]�
ǈ��e�[CF �D�q���vi��zF��ք�!Y$�B{c2^�S ��V���+����I�㼩j�rx�)q�L"�B�)�/S���Z���l�%`�&g�+�ci��^Sęik�l��]g[���q\TK�߮�Uje���:�-�2m�lV�%��j�q���P��%�l�-��za��s�U#�?��#$+��]OgI%)H��>+˖.���k�zC���^v�c%�m�;��Ĭfg�����ǃ�:o$џ�l��jr����}"G�j���ї��gP��2��vh¸U\S\,�
�>�X���&�k���Z�=���������_ N_q���T|��$l�Yq��=�h��%(���:fo@��8F��,��-�}9}G�;���F�נ5��k,Z�z��[KX����S�9��Q�-WQ�$�z�H5�q��:�������S������~�?����8�"�%��J>�R�2J�+UL����Ɠ�p���
�ї��9�k��>��PI���ܰ̏`6����J�%w���8���[��yݑ�Y����<E�E�^ؘ0�gx��r�Q���\��>������PG�)	��RN�ɰ�������,Ј�[y��=�Yv�Z���i	��Ȣ}u�i+���hD�93�
�>��{xp(�!�
Rk~�ڗGS�*������J�����T!W��Û�ic��Pu�b_x��U��&0Xܳ���*�(V	]���Y0c�	����8���nx�i�2]um��-�!f�Ճ`p塘f��h֋�����Uh�\+u��ƅ�2�L>^�!~A�(�&`ly*j�_l'�CS�\Vj��[?ӋZ\	�ڐ.��3ģL��؇�A��c�+�y!=�����Er9�ra����O"���Z����n��(Br2�gޗr6�Pȸ���e���*�q_[C�9e���RW�%�N�!^��rS��e�|���AΤ�?я_wn�|�c��xN�IV�䱗u0O���Ǩl���q�7��	�f��q�N�VQ�����U��C�$�c|h��5J�cQ���y��WW�Q�[ ���˽�qNW��ăy���Z�%$�Wy<UW0k1������M����1�*�ͼ?�1p�x���I+D��q*���FB�f�	R��[c@�D�_���"���P|�3�-eW��ĮV@��`�I��^;��ך�h8k��o�YGSĐyt_�c��Ȫ�K[?e�
���ᓣ��V��s��S�p�Dy��I�V(�U��]'�՝賠��c(D)g�ĎEƐ����*�_�ubq��h��!g��~�U���9��X��y0�N�=�N$����9_���d<ɲW���/j�X��ɻ����Ϗ'��^���I���7H�+Y��������H�)v�/X�z�Q�A>K�����G9	��ov��m_��Hz;d�\�lh�?��+�*���-�������M�pZm�M4B&�I7K{:�P�>�S�
qj*��HrT�3b��H?�\No�`���s�p��HyyTp4Rɴ`_�����%7�oy��j8�g'���5u14�';���G맥S��ڮ�Y�H��*􁜺w��pE�.���f�ED�S��PA����7i7�v�i���{E�qH�>�,/�ZNB�`<E��˱��6���zը>gr��PH�qb=���J[�G0�]ip�-�>g	���¯�$i�'� �泫��\�G�$a�*U�i�ȑHWertՂ�"�+%� ������w�籞��}��w�����j��v��@�(���Q�z}��2�d ��b��#'����`Y�K|?R�:CًR����)�l���b�j����	�"`�����:��.�ړ��r���4?׆4�(*t���|�/��0Ũ��M���B6��:%}�M�x�-u�uɺl�)~�8�j%�a��Bd<���`��G��,e���O����%7w������)�X�4����w�t��my���.�6NP���P,e�d2���ң +�j�_z�����§�rOZ��B^:]#o�Urܳ�f�bh���yk>���2�����un�X�<Gof����.�|l!K0�~iAc��j�N�0CʲA��-.e�(6�L{[ڏlw�9��\��7�]�(��gHmuO|,��>>@�J�� se��LN歝J1F0�;����	k������������h��g���F��fl�%qk ###��|�X" 3�W�g���; �6��ۼ��״�A$ӗ�h�蘀�=�5��@t���;l�� z���l
�T����������6%ᷧ�X����#�*^�-���w���AD���X�y�STtpOZ��TX�T��+1��E`1q<?��,��i��Y�'��1��"=V� Q�)��T���j�<��u-]\�K�ôD��A��_��� J�\	,E��=yR��r�U�I4P՝�"F��GJ���P�8�5�8e���G����1�A/�������Ze ����cdٛ�ߠ�w�L�Ao~u�v4�Z�;�K5�FT�Z�ڕ��z56�uu�O��;�������ħ����i��t)1�_	�W��?�k���ԭ׎�~�J<q�
C��R��I���H�����MAԥ���@P�� zH�:j�8��m� P�MO� C=��̇%Ɏ?��n�+��j��P���u�c�9jL�0����C[~}8
�cg����:����dPY����E7���F/��'�/���Qho�i|��i�����a\Y��^L���I=���"e62��FNN��?H.�� �s��'�qh,��#�������C�����8C���V�2����Ǩ�s��)zza�z5$*��T�m���z������@��YF��
�N��Çh�^�MNW�;Q֚=����բ|Ø}�5jF���7�0� �kC/5���#(V�lS��#m�F�H��,��|���: V�CX����t�x=חPT�_>�,j8���L�o<�+��hm��oL��f	bvy�eC�7��z�����%_����jI	��	�p8f'&|���m�I�'^耞Ɖ!��vMU��D�!4����E3b؛��Q�I