��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F��������n�BJ�F���U�FW9d����T�+�wt3��^��r�q;\��af�י,��9NL���ٴ�[�Z��^��Jy���0�T����l|�x�5#B�o* ��J/�CO������|�)6b,P;����t��ew�u��5�v�u�E�8����R�oIk�����Wb�A1���5��r�5Hڜ �r�n+��MS5��n��þ�|R1��������E�%��0E���;%�6�׸ۈ�6��:�!�#��L�jT�a�S�N�LS�[�&Ϫ���]/��nm� 8K� 7�H�be��
@��1>��?���X�U��&��P4
��J��tz�6�^�O�A��S�������EjS�V�6�$�g)�H!�uA�����.����c:k���:J�G�y�*aio������6M�pʫ��QZkw5~��ΰ <�z���i����Y�T�w-�q$��k�d�V�5i��[�r6t�`?�.�^�v�
��l�;�y/��y6�]*T�۔"N��d�V۬����/S[�B�U��7 a��p~q������~�5�LPؐ�V�T��?*�ؓ�C�r�����	�].o������߽o8+\i+�`K��+darwEi�JI��4?�}͍�<<�,�j��'��u��K�C���=a�X̉��37�Z?�(ȣ�$��Yl\e���=~�Xa��s	 -~����w�N���,v-�xa��$a2��hA$]��g���[\�7�x���{�MO|���1Wc���C��e,m�"��$�O��
	��M_O�~���jCL�"����V��P�h�Jm�_E��HaT0CS��&�L1<LJ�ګg 9Tp���N�Hm�}r�NBa<��9����-L��s�/�ap6@^߇T��!�3��`�[�� [ݭ��O�>F��� ���&�	��A�A��.V�Sk^�%�M������P ���v׮���w��]���B��(�	�r>���a������{8��Q5��}�;�9k��,M,���=�}�h��W�)@�܎w�B���Kt��	 �b8�V������^o���M�O���D��$���.�x��L�\E��{���7�ȍ/�$,̌�nj`�(��]Ks[��[B��Y�-N[lnZu��%~���e���=()�8�(��(�
X%n�1�]����N5a<�=P	�[��ð�����y�|T:��4�ybe} U2�I�BG`7>q� "©�#o�V�t4h!�$Dw�L�Ȼ�4�"F��[A[��`��W�"&\�f�2��S���V��N���6��& o�W3�pZ�AGꇪ<���r7v�>c��p�dn�l��=P��� ��#��{L�5}��_�ޢ�NZ��/W{�,���������.�L@�Ǔ�2���!�1-Y�;]��?�|H��2���BKE�*�����Y���-M�\�8�� 8�fwt-�,�dQC�D��8���k
�l�O��6,5�z�<G�$J���~{pVr$~���
|��s%i2�	c�]����D���ޒ����OkѲ^3��3U�'�Dr���f�sw(�,�44��Q�x%Y��:VL�j+��+�O��.�"A3���'��+�� F8v�SW�-��UZ��R���������a?���NӀ.�&��^�L���ά	Y��]#�|�`!�����`��Q7���v�Qm��#4�b��R�O�/�X����_�G���T���=�Q�3O�Q�d�}A�Ѣ>Y�z�g`��p�XӠ1|zCE� �L@X����Vh�+bò����E���>"�m���k����~���腔(�y��1.(e�`��ؤ�J����6�?�g��$(�)H3���seG�&I�1�%�x��ʂ�+x�r76HV|H���2��Se��z���EQn��k1�I�=�hi�B�u����K���f�&�1X�U��b�A�%�f�ܕ�P%J��w�z�h��]٥Y���Ɏ@�����ߓ�}M��������
�[N~;⇖���+���[
"Je�x���x.M@Q�����\������IDa9��O~^p@�B��B+g���M������^�G	��O�-_b(�L�09i4�=�:���h�K�u"%��:k��@V� !��6���4��j�᷿?��:�M���Q����^���c�?+�o3&VB�Vj%j��1����n(ʰ��� w���~[�8c9�CY�3g���W�尲Ri/���$!�c|P��U-��p����8:y8��/-t�i��I��6r�ʴ�?<���{��Q����69�����rJ���}�Rɭ���-����|l�+)�3��S��o�`��
�z�~�C-��VƘ�\g�F��P���OW�`%��Ķ����a>��3Ǔr6��( � �[�is��!�&�5�ř,�5e�0�%�l
�ȥ����N�6
�u'u�524A�����4Ӱ������Ʋ$���{�Qe�"U�q�1� c�=�
c贈��?`8�����vBw���L®9~�7l����C��y�U��uF �mG/�<�z��RU���Jk�Z-r��tQDVǀ)�a,�"Q�j�#'B��G �p��RI��m]�#�61��v/}u�S[�+����C&�|������K��%����8�1
�7OVAm'[^qX�"�a�a�m��/|3�✞$�������d�+�V����=��W+��g��E�׉���I-r'v.3������N!z'���r%�"�j�n��ćs��r+��l�#�#��~�={d�m�r
���8�'�sEG)�"W��ҽp�8[�(�g�� �t����c�׹�w�ö�V[a�����<��N��>�
"�������r���� R4��j�O��'�X{&��댝�B�!�t���CJ~���,́�]r���T r	�ĚN��Ǟ�i�Ng� @P"e�C��|�5��Z1�K����J��V������?�o�j����c9F��щd�Tq݈�sW����#������50�g��pA��Rd�����*����~z��`����(�R��x�6H����]��l{O�x7��-E�!�� F�s������%���g�fVH�7\��wY#�F?5��<��"S���}��
|`+�t���ס`X# ��h��pߧ_\��B�����D	bp�18�r�c�F�e�� �*a7�sc2D�c�X�0E
i���DU%J�Ɉ�?�2�����Tk�߃=]3��ۄ��/���W�_:�AM"M��"���t�m�(t�����$����IIO�Sh