��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�y�L�-��T��{�-�md�}��M[�xЎ�Y�^�JS�ڣ�mYlY�����n��B�}@�u�н�~�s������r��FA�%E�����������DJ
?�G�%�	��0��O�N�O��0Gy%>'���P^Id@x0)@^(��#
k�]5e���9XCN)��+�
�z0�d���E�e8��Pa��*=b�ਊX\n�h�T�y�Hy�qK��	���WT��,�/Ju0i5+����[�Ym+nUl- e]�z?;��+/��׫d0I���6!�q���4������-��d�� XP��'�/٪���1�@v������#L�~c\"�V_ȸ뚥�N��C������ْJsh"�Ln��v<+�a�� Y���Ҷ(���ތwb����U���ey�
6���&Q��\�&!O̸h��B��uig�`		�J>�Ԣ�h?R-�N� ���J�v_����Fq���r����􂼙ޱo��I�|�:�r3/W��!�����2d pt"s��$r/&e��. �\S����J�v٘r̻U�azp��H>(��Bv���Gh�s�a{U�*Wy	Y�U�]S�,(uUJ���>������J4���S�p��줉����_l�����K�1��첽@��Ve���.=���ʚx0�_���| � ��i'�%o.�WP�QbSoZԷ7�zY�~�G_kڞI�(�)N��N��ŘŃ�W�I%^���
�"�T� -�ȴX��%�(�ҙ�7����fd��ͭb�2�*��`M���P�Uw�n+�Nj[���C2	)2.H�i�F@b���{�}I�Mq~h���Ҥs��V���Д�����.*��H�T{o�8��McQT2���?���������8��ٞ=Tĺ�)PI/��1m� �l���L�8e���:��R��I�5'�X���K�:�wYf1��STݔ�I�z�A��fp��kiZ���J�Q�u}1��XBj 微������C_O�bMh�)����݌V�՘�����2�(�jS�l�%r�k"�KE $)ajY2 &���r*�����(�y0��d��R���1�<,F::y�ݛE�W�"�}{j�	HS'�M�Q�-	���P���]y����/+#��]����_�SN���?A}%�I��H������f�T� ��9�`N��y1��Bۇ��㦑��$���ؘw9a�3K�7ޅ�j[��e�V(Rg3��wf��B/�?�n��ʺ>��MmF	U�&��,��&�%a7��*U�b���6��G�SP�ޗ���՞-q�\f��=)� ��5����)��D����*��I3��T��M&�\��3h�Hb�/D`P����bU���s�����+��X���}�Q����dzkRl�(5�ސ�`?r3�t�]i�~YDvci��:b��m�Z9�O�p�y�Y0u���4��6���K�ո=l6\�c�l�ȩ�lwXk����B,r��������/�^�������1;���!��tun���FX�Is�/���l��4,IDIP�.)h��8`�B/p�˷e�%��3X�� Hgv��s D%�4��_�/�y���h�;3ޟ���z�� ���e���l2��(.�|BR�Zb��ࡺ�33Et5'�q��2�[�E˛��F���N]�k�lf�R #��{o���d��GU��iݐ*�h��W��ud@����^x���w[W�>�
�vh4/TSVCq�G{���&� ��4�b{��J��x�=��V��xB)��_����G.�6ǔ�����n%N����&."�����9�+~�V�7'�^.(��ϩ3��߮"�� T��m�ĤC��7�
L��59��[��J���O�&�\;wA�� ��}�2^�J��6+�{!=���đZ��&��-A�C9��9Ǥ;��.��[L���	��ȁ����w}k�F��G4��`�"0�U}G��I>��g��߽�8:$Tѝ���b6�����Vm����:ɠ�Hq�2��~D 鉯���P$yL�+��jpH�=w���6��44k����r�s9(�z�p�4 �y��}�� ɭ8���^k9�tE!c��|{��wE�:��}2%J���2�L��)��lwi[�iF��F�x3�.ţDf�-p�1aF��N[��?E4Ϻ����3��㇠Ӟz�B$iA��
��'�Us<Q�7��:-?�������p&��Jlüܴ�`&o ���u�Rܟ[{.Wҟ�����|�6�=d��	d�7�����W��p�L=�j=�����+����>{l��v�Q��X�#��A)�g�
�H(|����N;7Fe�"�^�Fhγr�T�'gب'J��w�Dmm�L�6��ׯE*f#;gl�
����4��^(��$�Ԩ6֜$<MW;9B\��R��c'^��O�y�=l�0r�7D������t����+$̈́�	-Q�����:�
�,�aD�z��]Jg�s�XیઙEy�VP�	��1ZGĎ���紶-Gn������ۙ��[:ίqfD��Ϳ�~�W��Ns�"oTo�lS�[���-����q7�ZT�$I*�S�Y�+R���j)�ռս4>��/̛�cy3�Op�yՆ~�o�\��@,ml�A�,q]$-�$�4����z����b���h�����#"�D�'�t`���A���}#��?��bӃ��F_�eс���!X̐s(ǛP�O(;E0Z<7��j�^�5,9����r�Ux�Ph9����+���֯{bӮȡ>�֙Ĝ78�tZ{�΄3��i�kj=�%�T�5PPl�6�;��S���]�̘S�����DJ��yH��K�]dP߃j��yssJ�e���P�H����q����W(HHɇ���Fd�`�{�_�/��c�dK��N�e߄J�ָc#yUi�+	��+6~ef��ۥ��F�qp)V�!�
�#�#пg��͹V��fߠö�!�g����4O݃�N@|�;k]` 	�i�b]tQ9F�Gg�� �8�<�̘���B�1,�,	X[�c��	qq��H��İK�%�lGe�
EE���B�I�~nғ[�����z2�S��6-9�!�r�.���"�=����@����� ק��H���G\R��i=ǴP��\%P����<�iW��Y�*�B��َM�=�T]c��x�H8��"Oq�۲���24����y�\�-��u���aI��h��ޅ۬h/X�k[�zz�����DEڷpWg B��8O���N%����������Q��.��������e
�ڹ����3�ώ&}����T�̽ �r���4��b�3���&H����T1��Վ���}54l���_��'�	��r�k]j��?�WI�c�[�l��:3����zs�
���V�s�*����:m��@@�r�	%�x��X���'I�&T��b�G��E]W���	� 9Ӿ���6��t@�t��d���4��~{���-۱���������D�o����G}���t���^t5��k%N�W�Ǵ��e5ԕ׸�3���K;�����x@w��R��$�'Ĺ3|��Y��9z�z�J62�(�����[K�zl0Ò�,��@����-������!T���m$���0��<&vƐ�B:\�S��~�}Ч�9�8E�8g��h��(�ZQr[�:n��'���$փc/"�k8�>���k+>�ڶ�s�W�"�!�i�|�f�:-�E�<6���Ăq��|�}ш�T(ΐHЌ[5�Og�����A�N$XKZI��?`B<8/�Rnx��[a)���9�'���)�nq\a�!n� ���/<M�4��,��H�a�K{��&�ҏˠ���w�Q�i��Ryw��,�Ćl�?R;�خ�`𳼐q����u�[���8_Gh�]��{^��J�j�*��.2�.cvh�b4�2��;j\��+|v���lR�i�U�e�0f��R���n�y�a��P��u�Vʋx�p�73j��Gz΅:��,2okF���9�� /�J��&���q>/0˂�5dw��Nt܇�����#\wƩ�Rn�����5ܰ��*:�5�#O'V��:���1�-��G�K*ΰ�Kt[�=}nM�c��j��?�Dh{�U��>��<G묊�K���d3gIŸXs�غjk5���;V6�@mAv�MG2Е�R8g�šoa��G��O�Y�b�(�eP�L�d�mU�C�.�4�\9f9����܇a�^W�	��dm��¾�ۦE���
�+���Y~:%�u;i�5}?H��q��[�t<�����O͇x��fng6Q�v��{
S��$Y�5����D�7��"׫O#h~3�1W`w�N�����;�y�W��m�@��B����c:I؉ߍåҨ��
�����b)������]�Jq��r 88Zn�a�ݏ�ZWX޾�����zo+�i�k�߬_���?�W�E�9�
�|�U���_WG�1B�����i���~�]徊��pgʑ�-}p�c��ܔ��D����`jP�.z�og����u��"������6s��:��N+�) ��6����Ǹ��׹��NH�z9���Q���� 0�N���9 ՐqT�"u���>_!2=>P��2u��`��7��� ��]W(����8l����_T���shv
���Ii�����?��v�s�G�N���F}�
zF@�r�������������Is/�Ȕ%kc�ٓ�$�^}���[tu�M<��oQ�\�Ҁ���D��Y��jM>D��a���0��-|��4�������'��d��Ep�o�� ݠ`�b��\BEr!~�	t�kXܚ��`��xr����_Tr��N��p]!���:e�Wz\dK��F��w��p���r�c�����Y`�ݮ���u���x�m��|�]��*U��4;�jC�ٛ�߃}W�>x�6 ���\���ۍ��� �D:���+��_J��O��2�`CMX�\A|�	˿+E�T�{-�hQ�#g3�G���E*�E �[Җԑ��3��k6D���M�C�+��h�]�&W� ]�e
,A�g�&���&drh��;���l���إ;ӠA"��/8hG�`M����x\\Q�Q�b���e�����1ȕ��PrD��Z��a�L q��S���J�?J6sh��K<���2�U��m�
[E8���I ���Ǔ����O̜~u�]��#��H��-54�ׂ� �j��&���)Jy���� .�>~u��;Ohk?��-
��jwѣi�y���u��2`���� �;�|�����I�/ӄR����\�#le(��$����2[!��5��l��=:�U��5O�?[�
��	�R]n�ӆ8�|�����Vlk;J~�"�*��(���X�7kV����^�δ,0T\�Kn��C'ވڶ�
��ȥ��>�MVQ�g�y�6�rټ���x"�c���8��v�ٵ�AO�>��.t!�-�@�iF��T0���Dl�SP2齇ǯ�Nr�	b���P�Z(8�p��MhmQ ͷ���ɑMz:��lEڦ��y�A���Љr�A8�q�V�O�O�/,��e2�:@�K#�W1[��`���l�a��
�+RK�(����S&C��ތ3���7ZG�Q�~ȷ3�SzI�6"/ڨ.�\�L�9���^�v�5���R��Q�d�V�|.\�����G��F_�{!��	W�GO*�kp�.���5b|�څAH�H�\ć�;Pt��ǃ|�#���HH��̻��;�����	�0q2j�g��w�YY�l7�D�I�r~|���7�̩3���j�����n[* ��/�<�����ǐH9P����*<�����n�^�4U�������}��cJ}sU����ggW@�.��X��2R��r�sZ��������2�{UoT��s+y�����IDJˣ�(m����M��Rް��z�X���)/��cg%�9����f{���X)m.��l�(J��� �$u@3�ZH���U�W-�!&��UY�$繍<�n���'��"��7��_hW�Q���q��>�N���7�9�_��Ё[��%D�U��*i$\x��6]|�)�648���m��,��Y	+�;p?��!a�:��a�A����/�O)Yp��l=�l����R����:�r�&¶ݔ��JH<�l��i H	�6չ 4����� @=g�*!4b���`��IV��ϟ��5I��Oi���>�������BEB(�!���X?��gZnk�4��1�L�� e�Yݏܿ��!�G�- �]1���Cb=�NLn��4��R@S6L���v����r1��:�C��w�+�r�a~fq�h�K��� $���@�^�?L�8��}=�N��x�8#Z�a��#�&9S���D�DG��om���g�P�W`T'�kh�����j3�]_���.̜��Yq7r�y���:�
ء�K�� ��Ɖ`��D��P�����D�1<�>��� d�̶�������jM��W� �"W&hg�+�����3C� �عؿ�*<��6>���ѯ��fЦ*��]l��e���?��$���S:�;�.tp���@����zi��\�"b�A�}s�X�r?*�ˬ'�Vuv)p_�}�	��%���ax�
)��ڙ�m[3(ث)�l\�V�LS�fb�0�����^8��!������L�.a
�g-`�G���%D���	h�d"��5M$�]�~^�y�	�U�Λ��1�	6>E-6≳�cr*]�d���=i��x���w�V�B���۞t3�j�����)c0kK<nF��8�b�/�-��m��f�����)j��jX�v#[7wz��镸5�7��V}3�]>F���y���X ��n���N���D�栲dx>�;x���[ߟϤ,텍�������[���yk��K�_�o񏛒@�I��IDNȗdN?X�¿A��z��[��D8��ՙ�{���wg:7�S�*���5�s�Ӫ�1ŀo"�n���aa)|������B��\:Oh�&�����{��ڴ�/����]�Km|��f"N�ㅨ���2%*�m
��x�wRF1�C�:�l�Z?��&�l��C����϶&�6����/]T��4a�p�c���]�z3��YSx��4*�[`��l��!^�Dmgqߘ
,���Cg4t��w�%�@�_�0>Ga��@�"R��h���8f!��J���O�2+�=�T�.�Ѵ"י�7�^�����q#	W�^۫_�Tϴ�h�� �k����>�O��;�z�]���|�P�駹�&�lN���B�'eJ�c��l�p��Ě���O�DN�Q�%Y�Ba YWύ��<9�6�8�O�3��l����D��Pnl�89:�/�PjA��/Q��w�c�U�7׿F�7�%e�������Ku����(�o�Q�M�0'�a�N|��X�-���}��?�:��ô�&�LW�S��,��GH0�vk?(+�Y�eY���:�b��E�����]�*�W�y�������h�pv� ��U1��Л��M�����a
�D��\ͅdKK�<Ys0���z�c��k>�\�$@����0��S���{�b�	�����R(�m*�{L��Q��io! ��{�M[���	�M�C7�K} �D�yD��1!zǀϳ�]b�le4�I�&�!�@�>�dt�P�;�9����r��$���]DQ;t�fJ=q�,7+\3������q������=�NT�ES�f8	�E��C��
�L�5Ͷdy>��_���+1��W���(�d̯.�ϳ{��[�⎑�rP���ϯq9{�lW?��������I��P͉��k 
���+}��j��Ħ����1���Ї���r`��iF��^�N˻v�,H�{(S+[��9!)l	;��VׇM%�/�5l�(�H�xENxd,����R}ja��8,�U5���ǚ�**)2`i�#̪�U�ϊ�n����!�So�Sm�������ya��]��������O:���������+>B�`�$ɍys׼���T����4��o�k�� !_�72l��>��2ZϿ�v붞V�+��6��l:�B�Uc���GS0f�em v��H����;i��~h�����Z!/�L��G���/�;Նۑt._tzJ���q�e�َ����� �=���$���H��-jpF���l2ܴT�����u���%��4}���q�v������z�i�����-�J��_�Z(����<�6n���40M����kVq�.����C�����/[nr,%���2�����[���O�y��)Y�
�wV����0��h����sh����(��Zo-R��C��'9�w�'p��xyȶ���]7s���F�Ǎh"����u�&Df�y���o��E[�5T�I����� m����� ����?r��_R��n���|z�ٸ�����쩧����}(A�v�l9�V�(u�o�F�Y�H�,Hq��Х�Y#nj�4h+K|��>�y��_�`fｔ!p꣒�֊#����L<e�Xt�������֑]hì�v�b�G�rY.���*T��k*�z��؊"!Z�%Q�H���*hF!�$�;�m��zk�~�j�#hݨ:4�zN��G�TQ:���N_������4��;
����|i�F-��X{;���L���q˟2�T���t��S z0��+��bd����u�������*���02��*r�������
�h&�d��V�����m�E��@@�L���'�5��{E�2�#�C�%bxSa���r_9Z��"�"izU�[���[[a�������v�L#�ˌDr��NP���[v�+Peo�t�)�h��D���r1�UR'���:��%n�8y��{S}���Iq��O�y6#K�A��wq:�i����,��9���`�����SJ67�~�N�Rд��� *I|�b��e�'s$����a��/V^C�L��ai�G5��#�K�?��ț/t"Ȓdγ�D6��P��c5�,<+D�{v�^Li�WbX���T��"º��V���)N���_����L���u]�x�'US�4vYA<fļ_���rG�����o�>y�=W�� �y~�%��*���:�xoC)���9���ɰ�\��,걞�0E�F'o�%���5�u1��eFz�ލ��vLXm��ۡZ$ٹP*qCy��,o0�A�9�k�Ӵ�Z؝�w�>�/<�>@��5��w��[�n*L��+��ٚ��kKrf���h<��EO}Zk�t	*�֍���9�q��鍦L����;��j
F�V�O�y�'�^2߈���h��j�D��Դ<� RD�7v���ս9h. �����ZU��jP 1C�=
�̳�:�nP超�������������jΗ$����?�"/�����g��6��pjp<���ُ���%�:YE�bT	�����Z��.��3��:��\�q�-*h��N�ǊCկъ{�R8V8l�nԝ���-�v�B�URd�[U�%�TnW1_���"��԰z��m�72�¢�w�;Y#�	��K�[HI��M5H��!s�=I�;�W%�^��BKCݥ��s��r�'�1����hN�
�K�F�39\2?B� ��P
`H��D:=A`d�>�t��TV�t��@3�ǡ���~��sncsO�6�nBc�m<F߮���p��1�bD`���Q�[kE\�#y[|��-x�r����ϓ�ERw�x�l�c���y��+�C��4T��H�h@�y[��[%3��Ȏ�]g1���Ǟq���s��Wq�"�r� ����`��V9]�b)�߁�,�0��ak��z�Gƨ���G|о)������6i_�@��ϩP���L�ZlN��mY�<��w�bq����%�w��Du8H.a�#�տCg��va����=5Ϋ�/��� Nu8��Q���Ҥg���	�x)��x[��'�cC\noL�NZ}��1?�š�ܶė�L)�9��ɚ�>���>����)r������"e� ��L���	pv3�K4�f�s0���'޸j��W_~)W~�[^v�s�����ko��CK��©X��@<�,Ru��@�-�d����s�=����0��ا�e2w;�Pe���:I�5"1�@u�Y��AZ
�?�y�>yG�[bCx^̛��wfx������O��p�[?GP��G�����R�<�{n����EϿ�ʿ�0���VPU� = Pt:Tn����s�~eޣ�'��T��:��_�����%��Z�l���|��?�����o�v �ʋ�?Ʋ�B�����^��G\�
�:s�sN�*ˠ̬k��
�y&��# o>�����5�e&g`�)~����"�����{Q��&mR��������/��w}��N�c ��)���6q~$�,���r	��ID�l/ ���	b�~_��X�p��(7�s>jf�eW�P�7��5��혌��&B<��&5����\W�o��{��h�E�7��jVj�Tv�|L�{��p<����2�+U��ž_�jr,�)6n�J��|uɥ�i^��X,��)�Eq�m��m����8h(;�7C<h�:Ւdp �P�RU�/Xܕڙ�U��B�{I��Ǚ��O��7��?�y��]�L'f��Ê����BW�r�]�ɕ�<\�޷``�W���=&+8�A{���w3�<O)	���q��`�s]���N��r��V:��N�="�T��C+�>)�*���;��i��X�β�a�6��~�:-0���V햟4w\�yӓ�䍷ai��j�~藎��򲚾��/�%���X�)B�)�L��]�K[�	�� w{ҵ���7@�M���E�
��,?��Nf�r�7��eVQw|���э���I�A?)��m	�1��Ͼ�Z�v(��4/�A�(JF�ӮG��3 ����?��[D|½>Y΀�8�@��:�ڵ��hh��hzlX!J�H�9I�M��>������EpQ�<�8�[Sޘ��dnLa$Y����t��̓���M�����;F�9��<�䨒������j��P�bl1�v��0��_hV��*���S1�}ڥ7d@�U�)lnE/��ˈ��l1�:R՟;���m���1+J��s�8�����ۅk�/�x#E
͎j��>���(�����'|�9oG~�����C�FZ�O�Vk�Xuk��D��2�P��:�]4g)��dE��b��=��v��n��գ�<�͈�_�,}�W��Bjf�lOѱ H�ӁňE�C�l����/������t��'���e<�;G*ͰQi�#��_h�k�b��SSNȁ�w�"k�-�t�q�����'�������1�����<WA��,�d�N��LhW������C����M�)���V5L�B��q����b�j��B-��u-3�W����c^�?n�)�?��a$�ı�"m�kٮߞ���;S2:?�¡�b�L-Z�Kڕ��9����M 8�DG�1��uC�[b�
��oל1���l,�}.6]�k��4z�PPPF����
Ε��2֘⻧�罒L�Y��2��0jvM��ڣS8�ī��%�Ƙ��2"�N��`0�����b@������q����WT�iƸ�	�%şP���\z	�m�w�T0�D�ٮ�M$5Q�C��	ѡ)�U�L��1�fV,��z#�W?�~����`���hJ�ݲƉS/����Ӄ�~���u?�y)`�K�]/̊��P���,ݣ�1ѣ~5��ě�	�ْ��k;�Ԓ�����d�IA��߂vD5�K�H�֫3N��R�ߕ������2-l���OB],��HL'h�*B���#�ur�w��oDJ_��F�,���Pdvw֚��bb��tOy�PPzu�`߼��% s뽼�/�5Qh�0�u�{wz$%�V[�Ͷ+�-˂�B�$�W�aHH�
D��f��j�z���VF�n\#!���jq��j�4�EG=!;�:���f�ѕ-�Sn bp��7�s�sL)���:�)�PЇ������+����p�7��@�Q��.�D<�m�ڝ��%/��ubn�زf��X�'�X�.׍�Y� �EI\CE$&���o���J}��}�$9�y��olJcs/��e�x;	T ��ڞT�ʘZА�;aR�lX�x�t��jC��
�v�S"{��R�b��l}q2�)�B���#�^���M;�Z�3ed�Рɹ�2T5�h&f|;hP7]5<�̑�3/��1�?�<{���A��h/��::�F����93�w$U=c�������m8�����J��e�,f�4~�B��_���x/���SN���ۓ��+綣!�v�QM7��q)r\F����#X���T*1�%,��u�*z��C�`��D�=Ż���H� �Y��\�>�s[�Y-�@Kti{��+4�x�J)�<��\�S����� �ȟ.\�~4�rGݢ�p��f������m����Ok��M#EK�@)��tZ
B���l�:@~�Z�)Rn��YS�,6]�#ߊ� �T�x�<�X4��Þ��:�#�����
����,���LA��}��r>���,#D⠼���Ύ�`	�@����JK��!�p��?Ww�m;��k8�������/B/3�E���}�88'\m0aM�3$��t��pPU+h:a'��ҐVz�]��pV��)u��� �d!����>�8�'9d&LS[� >�x^��O<2����=��ﹾ�B�����N,�k�g�9��d.M�� (���`����0�%:�x����%��&}if���s� ""������m�����x�3���~�7-[��q��e7ulE����ю���_6荡�j��� WUG瑵�}sd��$���S�K�΋f�ǥOIWw{��?�>�xX�O ��E�݊�$��`i�,��ͫBOׁ�z��~7�`vϙv�9��=dW"3�I-������<�j���]�7E�;�ϸ���f�f2 )?��l���J�_�Zi���Pa����~�+D!g�p"}�Q���j��D�PpV~X�b��&��s�QtӪF�R�@���z�F/A��o(w�l8o�hz����NwNm�Y9K�@�����"d�d�/M����5������`�B������^L�m�9}�������M��T*i�BW��k$�a�U#�#���؋as�"sj"��31��s.��m��=4�5چ���(��O�"��n��c��ג1�l/V���̙o�V��!:���2�Q�����5�G3�+��N�܃�p�.���~�$H�<z%���*�!v��]?�خ�i|M�Q��P<0�B?�
��:�v�y�F}Z�9�Z:d�,ȯ(��*$+i���q?���vש�}�t�#�$����5�O���	5��ǯ���4j0�R8Riϐ���>���,.Wv����|��e4@uN��->�k�̊�?ݕ��
F�Kl�Ѯ��K�sY�-`����(`3��M�t��Ӗ�fǝ-ϝJ�����D�Z#�c���c{�����L�3����^n����C�lXo,�hwG���m���e��ӊ�BDYōj���]sD���/��ɠ:kYe�C�ꕁ:���XF<�d�~�Z�v�UkU��p�2ͽ
�$?�p�y�"[�E+�J>Uۥ�_׽�W�����:��x�j�)���G�����0���3�7�C�ֱ�,�*"wG"���S��n�)!�]��&�~�@Z��5���gзV�f��טo�;�����MT �k]_���c�D��)c�C|(�Zi��
=�Sk�W�F׼Gu@Ә�)S����]-��F������ʉ����#��Ě�[���u4q�V��m�O��A��$�QBՖ.��¬�%�F�D0�����Q[��K�d`az�:^�4v���mT�g�M�fO ��^8�;)��K{�O�uM�_O�s1�] ��r7k�ܩS)5_��)8#e�Ψ^fUU~ϐ�жd-Z�tU��M��%�R�r��̇��R����S��� ��m�b�s#�/�[#.�b�L�G��<�����q�����`}�x&\�i�g�������5�LR�b2��e]2�[8�ʛ�c��������̴xrz��%-9x;���y_h�C�jA����N_��E����sbZ�B�m��@k�<	m��1�����90��k*�^ZX�7{8'W�|�#BV������
���M�f�П�@��/����)�|��w�$�,�po�D�C��!�W��Dj�V�N/T�U�?�`�'.K���^��f��Q�m����*�N8l�R��3�!�ʬ.3����8P��j_n�'k`���	ر�� b�[�fٙI?)Wo�Qr���e���/׌�� ��� ��U[<�lƅj'�VD9{XT	c���Ǯ��Pg�=��;Lp�cmh���"��d�{C������?���-��Y S��I�n�y��G��7��Z��u��Ak.���nE�>c�c��8���k@�x��W]�x�"�GD�>�Dar����z(��ܤC.�M���c-�L%���/S�o���	�L��G/{~����E����шQ�rѭl����L�e��2�7)�;O��]'pR�*���Đ(��EA�(��4X|>��%Cf�S��۪_u&*��Ӿ�W������gtԕ��w\����.�
��>ON}�`�ߞ�j��ݓ� ��dd*�할����0���,��jy��TٕM$�?f���ty�� �oA��6'#�|#r^��6	 b��܊��Ҋߒe�vj�����L��5虊"pS����t6������;���m�4����4�J�[�V����B�O������sN�i�Y׻�k
V��=��Y֙>r��a�K�A��U���cf:��@�$rm���6��))H�k�MZI��eW�Ę���B./΄�6��0��D�!�_���F��a�Y���C��Nn�!�a�����S�;��P��^���ui��L5����ۨ�#K��](r<�6�$�����e������ᔔ���94�5����M.�#�0���(%�W�C�==.��k/�[�ޖ��l�/����T�����&
����Q�zU*�)u[�l>{H��*̢O���t�G
� _e��|c��cꗀ�>wݞպ��sL�7�1���Ƀ�:n�Ѓ`iॣ����,��8����o�Q��M��ʀr����������L�G�%��+�N�x���x �l�P�v!�����Z��+�򧱰ijR �F��V�	��ѳ�����v�_��.�Hu���J'oH �'��jh�(����'w����2f���[{+�{�hjM��P��GA>�*0���� ��C��H)f`=��\������_�Ϸ_�;E9�Ԃ�:?����&��Ȅ2�?��xQm�ZI��n�v۷l_� =��1�MARF���,*o�����F=��v������������'2�G�wE�@�}���H������t�����M���'�'�"�{���nNr=��:pl�R�c��P����N���gd@�"c�퓀S+C1���'��!��wZ`��c<3/��?�_U�#b�)����h� 	نyK�u�r"�3�2���߬��un��g��k�͋���y������>��f�Н[MB~]~��ӝvd�P6��[O��߿U*fEa����|F����,�cJ�bȼ܍�Mn4��J����i>2���Vrhغk̝i2��<�ۍ��b2��%;�L������P#��H>���W�/���I�pPA��y�>,��χHK���m�ųɬ��E�]�"���L���sWf�G%pj:+ \>m��[#�H; R�~�,s�V�+)~�ԏ��%|k�� >�2��Ick��ᆇ�IE"�0�V���ż��5�^~�d�{1ͰB�s�F)��U2	ʐ �2��u�`�1͈7A��ED�S����c���ᤋC؝Iz�DH��΂0��>�1���m���F*����q�>����|��f[
�/�f�ʑ{�C�4�MG��'�q=�-⢒�ΤzI��-7���wu��l���Kp9kK�͖��!�ʬ2�5��������i����t��˪b����/�Ep��+R�<E��A��Ir�_���L�����5��� 23�h��VF�q�v:��c?���[1ᔐ�Ù���e������Nx�$�h���Dk(-��ݕ���T7��!�h�>M��j�fwɚ?�b�^Q/4%.��>K�>Р�a_�����؏��[a1!s�(�5X�Zs����c��BM�t3�MN��E� _g!b��<�^ `v���)AI��o�`f�����7�#�bR��`^�� ��m���oT���l1�(��/;$H�#u�4ƨ_`��$�Ґ����!9�^�/pa�F����V�4ܣ��J�v�Αh4���=�"��e�N�����\x4��O�5S�ߢQ��F����7 c��e��3�؆���vg��m�a%���?�繤H&ݜ'q�cP]J�_]j\'��+�ҁ��y�p�0Ų��D�Ԭ"�͍e
 ���Ы��̋�^K)8��I�X[d���
�j�P&�p}j����,25�^s�b����V�`J�N3��=�x�����Ƃ�hC/���<�of�����*VC%��hj�
��wF�Kf�/�a��t2L�b��ٖ�G<���W٧��Z��^��I�踸֌g��ȃ��.�\EbZ��+=q���A�5��s���+I7�Lhѥ��4vޓ��4Ey�vH�FU>�:1��?�����<�Y/����#�]PF��� ��>�x�O)G��9��d��W�A&��Cj��=!���3�vf�?�s`������BM