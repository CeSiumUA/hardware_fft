��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���=��;u�#��� hH����<�C�l�1��9��� ��;��*~�~� �B𨰹TPvd��w0����Bm�`�~:����&�������d�6�.�����&[�R&MK��MU �
V0mc*�9���v�kո�p���@?�+���O��p���U[��?,^!���0�^�E�CMY��&���7B)�P��f�ꅿ08��h�Zx�~�����O+���B�s��s��p [��#�{�2+d4u8�Hd���F9�C���Vi��6�̒�*�k+��׃"�a�}�\�KT���-"fsQdXt��C�������Ml�ۢv��3��;�����g�bD�7�<+�7�ۏ�\�i!�;����E�j�ƪ��x+^��5M��%+�������2���n	�R�K��=���n�	�)ZGt���N3�LM�b&4�I^��9Ȧee֍5H� @�����^���uy�+��NG)��)��������cP��ǫ��>C��\��e̀��F�aO�+J럂}����7�`��I�T-;.�3��L���"xM4�m��&Z�f�9.�^���-�P�[=���[��C�	���B	���a�*|`��Ʋ��qjɐ�?t?���˔�.؎� �cf.yd�`�gHyR�+ª�?|��JG�F���HNBW�yp��g�2����]k�q�Dɀu�ڧ��;���p����/u�����$�U�He�
�X@J���C��m
�5���~bח4H�N���Z~
�d�6�c(;�<���";��fJ�|�О0&#~A��f�|lp�[2���Y)%����;�Z?���%?	��{9��r=T�x^
�/���@@�]aN�?ۦ%��F�7%띗����`���d+W��\��۟b��DU��Pc�gA��^ߗ���O��p�De�<7/�t��to��D9�%�#��E��Vbz?#� 	IQ��B�I���Q���5ü�"�M�J�v�K&������
[H� ù(�D�;��s�6�*6b�=��������cwbKj�����%o}�d�G���UNL|XQK���4�.� �2��rџl�2��*l�A�����pl	F. %#�c'��&�zA�ͣ�m�.��$���Q���3�S��{msN6��� e��L8�p/2��R��M
X3֘���*���}�������{�2mE Y�/zm\���s�R�ح:A}�%��*��$��t�F1�V�������f�hA
���������mK�X��u/����Ȱ��0SЪ��TD�w�1�����ﰮ�!���D���u  �(�Gh�Ynbt��"U���ޖ�<N�2@�Z|��Q��.��&n.��i��"4�\�����	�v�p9G�IA�ʟ�?Z�ש�*	k��+v�>�P����Ƅ4�.%�+�]�=M��1\|E<-y�g��qd���䉼�d,���E$�`�W��gD�T�h"�^ۻn�k̩��ly}F塕W�B���?��m�j�b�P����Ou�]��p"��U���Q�l1V~\h&�'O�x,��/ˢ�e�Q�E؎(�Śt�� yaP�޹Mmv��c��W�j��MՋ�z�/:�2�r���=�&Z]�,�+�[�`\l�z�:��-���X1E`hd&���O��r/�Z8�}�| ��1�J��j����3��bSz4v�Hpt���22���k�147iC8սPl�X�o����GKA�Xʄ�e4uqj������L��ҧgޠ��HR(��E,L���c�����-�4?1���*Fª���z6���9��f�m@�_9f�fj����4X�s��=M��P
�4���}d@��� 435K�0m�o7ʙ�[~��ֶJ�q�w�۩�"A���N)�}��1lO�bP�&6��p�iq!�,��ISpjB�5�]�P������n��c|�E���AVd���-�ue��Ll�b4f��8�΀ѡ/��r�!����XJ��萅ZsLZ9��T�����i���ۊ�:#���S������	F�����Tӡ����-D��B���԰�N��˞�#�~?d�T���Ʈ���$�!~�K�q;�����&��˫(��$sgy�Z�"̻D�툻�`.�16�O��K������(}"�}�ԉ�&F�efo���/�����)��@?t�3���5�V�GF?�����p4*� ��6�z�*���P����E��F(H��~5����%�(�e:�:�Ks��@B�+��z�ʰ�
N����{��	rn�����&���KgL�I�=�!�(�+O^#WZ��25~&�V��5A}ĈtJ��:��Ǭ�k�̮)
ijZ���A�ʉԛ�o�^��&96D���	o����C�+��8��dQV ��Fը���H`��σpU�L�^��h�A�}�`IUn6�ֻ��� ��$�.�*tȮ#=s>BW��pvmq��82
�O�$wʖ����U��NG81b.s����3���2j����4�.�/0tsqnt����a�Xf>[����͊+%��UW&/��s^��c3�ȷ/�rۢ�Y��ħ��<�5����2�xae��J��sN]�S��+ř��f2�p��3+�[�6�~_b4�q�k��M�*�F�sԳ��R��6���:4��Z���IS���c����$P��QFe�������ܼ6�@ރ#%ǥX����%��6U��|�G�ڱ�����u��nW8�Ee��(��x'�ƙ�<�I4-���jcy9�z���@vq�:˙�
SH���,S� 鸁2+~��!L�w_�I5�����yO��X�b�t3��o*(��|s\+��;s��i?��~EY �l��U���ԫ�~<��oC�]j���	�ppH�B���;��v������~8N���%;��p9w��
����u���Y�㑑���Q��#��e����'��dXP>	�'�yn{��#B%7�¶В��Z�X��Tʠ�;���z�ll%�xA�.�+]�	�}tӭ���ޱ���������چ��k��RB�W88ƚC�Wm�S�m7X_歌Wm6c���$��U�\^�{g�����E ��&��5~;��(�P��p�j�����=�[�n�x���m��u���g�{�ѳ�j�+�À
�<�{�wK-h�Q9��BD��k'b������z�OQ�;uϭ�L��� ��?�2�B	�y`�`5bD���������+ �����IƑ^dK���B�K��MUx�P}��h_E���Q���4 I���\N�ߏ�@���o��4�z?�D��#�,����6�5u� ��Gv��Ì氥\��1� ��hW$��Zڤ�sȫ1,ͯ�mV1�-9�|3�J��wR�M�G���o.%P�r"�)�z������|�u�O�lL`;�/�T������9��9�eJl&Z�A\��Q��3@�z���
���eΜB逯G������^ ,ܘsݵ|��;|5}r�C=>��2d2�Г��4��[�"'0�k&-J>����>�u4���x'_>����BXo��u�qu2#+'��Wa�=���D���f�[�p��Y�����)Ymp4��M���]��Z�⣟�܁E�o���Ddz�����3��d��f�(1�K/�L#�[��q�Z��
�1����W�u�_�$9�W���+��X�jk�x��{�(UB�f�蹑��>�٭�E�H����S<W��c�0�Sm�-�=6M*��h�b��Pg�����*a��@Q�C�F{N[2zgKp���C놼`�B����aT|�8�O����U'���?YP��EۯyW�<�`���=$��N�j=`EH�DJ+%���Nv0�fh&DI/U�F�P\��p�>'�Nz �i�W�e$M������,���D�=�� nj_k*J��fC>Z����9۶*��#�Bp~����tx�5�~5~�Rvi|%���$L\����ߐ�:' g��y��4�@?�:B����O�ྊ�N�c׫8���%�e��1
k?aH�,�����j�hR�L�\�[��Lʏ���ݒ�W�/*����_q�ڿY�'/�i��f���G:%ʀL�_6��Ӣ�ۯ��h�Z�.+����՛�V�.�2H�t ��S�d���R������+����2��#������ �+��J��
�/�	3蟶'K�ή�BX��6�Y<�(d+qƐ��ФW6$#Y����Av��c�_��}xj����1B?�c{��4��=���R;|m�\�''z� �;��w-�k�Fz|����G����v�c�����n0�VM�\L%GYx޴��� ��Y� ��ˠ'�q�3&�u&�)���<�dj�&u�P7���8��^)K N�"~�HQ������hϯ\u�$��c�z0��+ۂ�B�^�=�ro�����JU�<�MÐ���� ��'`�ߨVo�S_��zO�@J����*�<��Sd^y�<]��b1� ����l�<3�̶�ޜ�G��OﲼN�M���y=�Z��]��v�aD����{�T}QO���#R��9�c��Z8O>q�Oay��Awh�X_���ik���D�)i�]����P_��|Bo,OV��\,D�����z�s���wB��������f��2��-ܚ�y݊�W����㍽2ݙ[�S��剆*���Qe ���7��tC^hy�zi�jq�{����xb��޽",h��#�%BuA�\�e�����C�MΗ<�C���EQ��:��d���_�}|/r.!���U�ﲲ��������6��3�[�g�ʔ��!��ݺ@$F��@��E��	gӾ+ -G�Cƈ,�3�?��y��/��T������'�����m�"ˎP��B��l�c��\�Vr�� Ih�I�`���@7}��H�+A�|_�
����?/SY�-m�6Nzׂp���-���0� _Ω��r#	Bd��q����_W/�p�ki��B�������*@:��q���+�x�ݠ����lb�'P���߰/N�f
"����x�ׁw{�l�yK�0��G�7��z�(��F��]��O����"��tv�lm}XZh�)�qn�-�p_�~]B�5$:�Y1����	��9yFV���ǣ%���m����	��B]��r���H��v�^�R�Ċ7Lh�g�w�� 퉜!Z���ni��K�*�D8U�;�,7`��mH��K�'n遉� (��8b���3�B/ j�KTY�Wl[7���m-��MG`	�K)#�Ќ������{���$�T�𥨵ߠ1e�E��^]"Iql����@�j�7bJ�-'L�3�3jw��l�z�Hc�\i ��� @� ��OMw��(���~�8S����0���_[	�Z}{cc��..��ERM7q{x���-��g-�d�RM��R����g(��&(�'���^<T��}l��+	�e��n#�@\~M�ľa$=�;���D�+�$�h���%��c 7��a�9����*z���(ʈ޵�Y=|��a�B�^5�9�����L�&�2��I-��͜Y�9dC��I�~��h^����==�\�����k�P!������y�N����4gV���S��� ��}U�G~t�v-H����MG*��5��R��ꠒ���02�Ę��G5#�k�3rq�q�n��@>^���ڒ;ۓ{�}��Y;3���L�!7���z5_�]��h}���C��c=�͚v|��5��o �Ǉ8�.x���E��'R�Ӵ���w_��/c����mlA|>L)�]2n��轤:*�m�anlѿ�R�u�.ݦ���M�s���㺁\�}��>a�x�}���r�3Z��s49�(�1�!�r�&������'4.�ӧr����i.����ի;;@�]�X� {�Wy84��X^(�{v���Mz�wkD��Fҿh$	:G���^Gm�̫�x+�L���6�5sk��sY�OU~�D��>V8�ߊa��N=������6���7�6����P�����$d�G��c�m:yl��l`�i����X+UH7=������o��]�Y�^ǐf�����y��P�W�?՛�=��5����y�V�.A���������� ]'��*�^��Q�}|�������jCV\f�f��.����[`%����Z�aR�*�.-�x��	i+�y��Z��9����-�A�����\KwI?��~�n��S$�c�jJ)�j��z4���WB�
��H5���N	!�h65�{P���Q��daaaN3o�w�b�@]�b��Q��'���G����+�����w����;7���� lj#RTRDf�m�L1]J��P��� ����M W�j��7�C�q[D��z.�#ı�xՍ�Ĝ��q�X�eF�ȒD�f�8ҳ�7�<��}��5�*9�O^����#�����7�����X�1f��gq����GѺl�zJ�C�U���6��/ɏ�x+��7�P��)�Q�t�"�@�p�x�#�HQ/1R��� ���^���>[@��<���u�;kk��H�����=w�f������h� vKU�3�1m�_���-���FM�=)��N�FE��m�!�`-+4�����Bs�����X��Mf�������F�{��Ü�*��9�`�=k�.�CHXL)��lo_���ZW��#!mTr�*�F�-�3�c"�����\�����)�s��2���s��_������+�֔��X?�}±���>9�-�$1�`�����D��p�[���U�d�0I6�O]8UG0��pL�[%�]�z��\�๨���AS='}�^h�K@u��D��"ăB�&�4s5-A��!���s�y�b
ָ�l�W����n)��h�����!8� �wW�L����C��.}�:C���}��Ğ�@Q��]o��dY�	��I6ACr�c�/x�ع�E!��c,��_yx2Z~�}h�n-b�#�z�6<��"�������\�\�ڲ��� ���؆'�,"���k����%�Ɗ�������MV��\����-?�p����J�ϵ<��mj���rV�]M0�WԵ����}'}�,KC���$e����-�rh&��rh��,��D�x�EtQ��OR�."�.	�"F����e����m��4��# ������vA�A���{ǆ�=~	�Ʉ�p<NnY���˫ο�&�8��}tq���<~��8�ǉ��U$�������.��w0��X����S#�N��IV�t	��:��[�Bj��秫�"�a��x�=���aoi+	�<<�ڛ��L���׊ѕJ\f��3�ZP�V�rA�'�A� ��PeP���->��ǘ5y&�L}w��y�tpoy�d��wc��-��OС��d���7)��}]\�˵�yV=��o��*w�W�"u�z��u)��/;3��2�uy=O��t��� ����6?���-�^�0�zN}����?|	�մq��T��Y����v�>E�*r�!E�Z�Gݫe��;�`��+�5�!K�5wIpT��W��ҊU��h�����i༄�%�,̄��1gt����Y@ݭ�s�6�8g�����j�x�}(	��K������!X0?2`�b��u8Y���M�ߍ�>�7��O������sq��n��>ڰ��0ԗ�>�o��f�z4v�b(l�l	`�At�4�bb^Q��N�����G#4�M9A����#oF����Tur�$��1,[�Y$��8
y'���h
�+��R���_�m�d�A~$/c���߀�]�\�-�4���F��X�/�w����徚W%�]����Ȩ+Va*p����E����}S�o��.����6!ygƴ*�ű9� �t�ڐ�������x_�>��f�(��<:*Zc�h~I���h���/я�d%���I�����Z\�_���nM#�25���c�`�a�����y�����Uf����ZwS�m�cȪ �Ԥ��.��/w ?"_��tnp�����iN���d̮��ҖQ��㖆W�.�Ir)�+�s�ZFYl)��>�^�U7�פ��Y��P�����G#&-9,�3�\�F�{|�J�T��+p��$Zǻ�Gv��&��r�[�Q�5����`����%�e0w��')���������d��	I��`u��l��&u2R�{FӐ���!ȩ�~�2c=-*�"�-��^.�n3xO��,k�~�ܸ���g�~c��RK��~��KN�WR�k��S�I�@i`*�ԀS��ӝ�h��n��41��5U���+��1>k��Zv}�*�A��\����������
��?22���.�Ö�����Cjs�gaE}Q����[�b�n���UbȌ�	�@H'�oR�e#�t4����kF�V�~���z��..���۞��E���Rx��gw%xw�?+S����8��,�,l*q�B4˄�6M �O��|�����Va<H��r�q~Yl�z�:/��B�.�Zi@�-��r�z���S�>^����j�R�@U�����(�X���)2�#G�
���7$ݔ	0.f�����9B���a� Q���{tȢbˋ۫kC��%�^>A����[�q�?E�<���J[�h�!��Bnl"�h	��R�xQ��D C$�� )$�k�����s�B��/B�s�PŒpi�AFnbQ�D�Q+N<����L#��!g�?p���r=��*I�.-8q4`�j-�悎,f�I� �5��0k^;��%)���.;;�5�JQ�>д+
	N���I,3�<�������j7S�"x_`֝���P_X*�F�#0{�qW��G�Z���i�=晵y&)��ޱ��Sъ`z[5M`k�ߛ����K79�,ٱ�Gx-h�@��B���:��.ۋ��ͪ&��&>�9|~c��.J65Iϱ���iVԢb��8��N��S���o��I������j=��Q�MeR��zٝ7�V0
�e��%"U��sJV(D��{��C�]NPyJ��F�}OZk���)��%��h�!����a��/��"߃�1G���DP���A��F!�R����yslN���52�"E?����W��n��b�߁k��h7�O���5$f�'Q��I�oe�5�[�������Ik��d�Y�6�QB���D�̤Y�w(��_m>�e���������5t����m9���4��X(����Lӯv�"V=�^J(M���r�0��)��m�|8���D|W|{�PY���N"_�!R9�e
�6�7��=�	`�@��k�. f��Hy9[S�R~Ӆ��e�ފ��ǥ�_J��l)�p�������A��ksh���W(57(�G!�N�ɒ�0���g`�=�y�m���b�2dz���6|z�~K�Q��rB�m3E[n��!�4"�/��W�[�WEv��т�}*�-ޖ�tU�a�-�>�g)�Q�������z��H���;���?vk�M>Y�B�.vwU�}`��#
�2�&'���E`�T�X�F_��"e�D�01[��
��@�y����n|L"��{:EC�T��\���س�+��ؾ1ʈ��&���<�)���`MY�F�Ba��	��͚�����BQ�q����t^q�a{��y
<��^��FA�����BSڣN}��Ŝ�$:7vH^�/&SaG����}A�.��z������ID�(቗N�^�<�?d�"i���!#�8�Л�Z5d%�"N��Y/ A�	uN�dSL�^O�4U�Vy}��eP����#���b����TN<4f/���[��4A(+��A��'an#��l7+��Zюe6�J��缂����=eՎ�K��K=�)ɭN�� ��Z˰���i�j?A}����3liL�i_�d(	�h�c���B��U�7I>��s('	�ۺ�1Xߴ�G��2�o2�'>[���EN����P�̓� $��!8�pW'GxE�m9'�qqu��}�#�DK�<B����m�3��)9x�*��82B֊�|��Y��mi��@�������-��� �5��ҤZx��ypO��T��c�-h
9���Ⱥ�xa�����n	��}���y@�?	�{�Tt��]��6��6�j!w����k�.�/n�i�����-�d$ڏ]� ���� ����u��v���2��*��K�s'�غ����A��G����y�(�g��ԺP��M�[��CU�B�~���O{M�z�Ѓ�ݭ�-��,ѝ�Y��o������5A?�:I��P_p�j+$[��}a&��=rk��*Q��z��K%��?�7r�n��PS�\��Xv�B�Ձ��r�'�L5{�Y�ʀRB�g�/�\���
R���U%\n�|N6/�w#=�5���?=��~;wLm	��Ca狁-a
ztg��{�g�B 3���]p�JE:�"�c)rBR���˶��=�����_A�\S�A�At2��O���+f��q����
�ל_�^���*-��[l3��"D$�7r�k[^*ܟ����~@F0�������y��E�@�XR=�xG�<�do�l�v����a�b-=�c�J��'�P�ۆ*`��{.��.�����_
Jty��]�<�=�MW�gn�����=+~T��co�I5�,���ŕ���=3One�	�=��c��W�a���;�������.� e&���E������l��%� }H�!Vc�"��w�m�+���Խ����B�{͈r(�A����N������YǠ`����;��W���z�w{F�I�.]��!�םN5����R�W�z�v)d��`ޡ�{��7%�ΠJ���+2�n�gA�C�)��;�L����7C�!�oȃ�ڀѦ���݄�7`��M�aǂ��X�*a����S�T���A�ō4��cL� �axu\�֭���)�KĠ֛�X*�LZp�Х��%-+�yc�ß���Q��r�-��g��9[`
᜞b��`֍��'��5��Y�&뜁���O~�G�)Ӡn$%����d$mA���ҧ �5Ѳ�;��ٷ�Lwd�W�����=Eb2߮;��%k��G�{߸��s�r�$ң��}Q�gմ5���� 5ODI�oDTf��Bb����v��V��F$��m���A��jMĕ���*�6S[���Y��a/0�@���i4ͨz���M�M4��X>��̬�x��2�QtZ��Fc�7m��������G�a�������R6#����E��*��,���V�i� �X�o�*�{�W�\��}�\K�%_r���wm��ͪ	���Hˬ�&5�G��U�Q'�Q~t-!�û�<��÷��
 
p����K��Y���kR�Ђ��S[�C�.C��gF���SaG��U���蓮1�ݫ����)�� �\Y�լ~��Ґ����:G)��`'�7�74{����0$�}:?m�Z��9�� u2�ֈ3Ӥ�dQ�1[. y+�Tw�B摆Y�Sq0���z�k�%C_����Qr�o�e(0�sW��ta|n˟fHU�N|1�${`�A�翜Sq��)pU�SW�u��%�e���#��Y
�l2��I��e��I<G��Ą�5�`�݈�Lj�����,����yf�f)瑦��2+?��/�W��}�D���(VDh1�.�*C��$��e�ˏP�
:%/��������f�rg�Նj�On@_��]i����N+ͧ�Cq1 Ho$ܙ���S�I�
�ᨎ�k�L�*V�.�Ia�+��62��U��H�^ع��x�����`��������]�`����s��x{@{�ggV�T�c�20_S0;��mٹ��B�KI'��d�SAb���צ��� _l\!8�:���֐p"O�7`��j%�v�Z�
�;��t'KH�BkC�_LJQ�	��X�'1�����9��#,�� �3�?5��t�������	�E�Q���Bd�C��6���tP�ӧV�h4q�C�<d��>1��X�iT����HCA���fP
Ѯ3z��,�\���D����<�.t�w��4�P0lC�����]���<�Y���pf<_,I	�
����33A�KhXN�4�?���qN��j��,��o@n�Á>� W��.41H�b��B���o���zpU�PTW�b�����)#�)o�lRͯ��7&�o8ЙA�Lז����2B��i�8Ab0s��0�'���4Wg��N/��B���� �p7�w�a	�nΖ�pD�!�7����t�<ۻW�����2��	8u��#N���]��9U�����k��d�}~+�grC׫u��g:�Z��,R��J�f���#��˨�y���8����cl��/�kc�Z�5S�����%�T܀g%��^�^b�0#bQ���k^p0���X��
L�.PX�@JB3��6����p��/d��e>Lv�O�����1%�6�O���җ�)G��>��4��?�P"���k�!�`������k�YҔ�{efn{=�#aP�}ۄ�Ƒ�8��GJ]G�%2�7Ք�4��8�J�� x�#`�YhnC7^T����݅S	��Eܗ�������:�eh=O��᯶}"��+gGWu�倌�z �2l:a9'X�G�7=�]������ySm�G��`FS}�)lP=0��bCI,��E�K���çQܻ���E�ő�{1W�P����h'L�P4�@(��;�%��� �h	Ŀ�B�nn�x?��	4�6��G7�h�'�)�J��f�2%e�z�}����O@mbvG��_�r��v�Q���X����z���G�N\��+R���J4:͕��̇��!��_�	�TV}+��� g.� ��u�a�����& Q�m������JƎNS��`�sU�hk�@�\nv�3L�����7��Ql����})���l��h���nk�H�tm�.��hl�n$�%�����y�YE�+����5�f��O+C�9�s�ŗ�tv�����W��}Cg=��i�,��u~J�N���{8���㈌:!T]��.��F�[x~�g@�xё���@��-��U��5`�Y5�L���b�j@M�`���ܾ
�U�����B�+,X	��9�W�ُ94��őb�[�����f5�C׏M9~��6��gı�t��-!Ây�WL]ձ ��$Q��>�7%�(�!�����G��
�D�����|J�BBfSN庰o(�[E;E�-��},"(��V����-�g�Z�XbDo��១?�L��V��;�d�5f\D�^pA��Nn��=�"���O�߰J|Å3���>�v EH�K*6��#�)���Gabj 1ꬭ���x�f�[ߨ�`���=S=�T��$9
�_��oo��1��v��~�m���A<I���e��䃱o�|0.�Zن��!��'MU��I*��a�u�*��S�1�������Dz:OM1�,ɴst)���P����n��,n��2G�)�5�D�o���x�L�m4<Q�og.�*��Z���R�:P��EQ�`��K܋%.f�_��H������ia���"׎��pꋿ���b���4���#��=쯔�yts�y4��ti]䅦)Z��B�:@� �WR��%x�?Y��f��ݍ7�-��q�Ѝt)����X^-���)P�oh�Z�>�ߍq��}l�-cSv뎹��S�o�Xc�)����l=/�t��n]�"�g��l�\���8�֬�d^,F7|��b�M#�g@�U�����i�W���It�0��+;p9m�! kͻ�Q\'�"9�ZC�7OZ�lsL�JvФXN�����5�*�T��L��(F��{��L�-S��x��͎�0ퟏ���Y��K��2 :T�(C*Jmu�(����$��g�/��P��Q�%��X �'���Y(�(���[�We�p��v�H���Kn�~Y�d)�eŸ#�N(�]���$�Q�& �����wT�)z�J=��V`�����H�����XEz�Rmi����[��damT�#x&;X��"�W �pXY��̾������^�:�P�"�i)��X�A۳~�Rh���C�����m����R0^��(�ʦ���s]����IW1�K�Ob�F�-�0�:���f��`G~0���*�1p}�C��/w9>�_��b�ը�@|��ݔ�|��"���o]U�XǠu����.�q"J�f��=�j��	���5���[��by)I�w�j���r�Q��UJI�aM��b2.�Y�O^,�לC�/eL�x��u�|�$y{�bx��{K3_�t$�͚Q´e:�ck�5C�ˑ��XlmirUV�������+�xt�Č��se�xA���i� ��2D�� g��P]�ה��E�xv:�
��ZUk*���u���4�d�Ξ���݌�X�W�	i��ܷ�E�\w	����H��W�P'NeU!u��0�x���X�P�z~�a01���.��gk�{M[*�[*˪]�Y;�a��%����K���A�f�j����)V{3���zWw���l��ra�1;�!���n;���0����_L�����t;��9��bh^Nj�-��~�K)�@����^��6�����H\��R����>;�^���g��f�lFD��5�	��~mpDӉ]|�����0}�?�
�r��Ht�Q|��Miw7�$�<�T1��G%�vJSJ/Q�*y{KS+�� ��5���^g�v�v\<�ĴR\�k7"ⲏ�Sgu�����6�4j��`y��`n�\�����7��d/�u��wI�	�����H�u���'2�� N�wI?�!<s��w��vn�s�A��歷����֙�r�^`븬��&�p˳i'|��t���V5� ����GI9�:̑VC�n��2%�$����8%s`7�o���Rڤ�{�*p���"x.T�����	n���j�U����yNF��%
�e���۔̒LJ+p��6 ӯ��a�_��*�A�:<�;�d�@l�C#�I���O��d@�Ә��$��T��d���dEA^T4I���g�w2J��
ĩ0���ʅ�C1�r�tgU�?jR,�Tzz�q9����V�����lUj�����)�b�j�6yZ�����='^ �}%��Yb���\��q���X�.oKKj�4��Dk����~��Ң��'���S�����B��,�*˵&͈��<�T꒪^]��*e�z!|ga��<\�X���:\�/v�*l��he[�J���"!�h�-��'l?f��}�TE����S���{���c"��@���i�y�{�v�y��qPEg]K���HPSN`X���f�9�����)��v�I� �3lM'Nn̨�֣5�j�p��u�"��f٤e;%����\��q�72�^�G/�E1-Bْ��keeQ��G�ugޣ�_��-G!�M1C��؜p���C�w�@Gb�k�vb�J�r�?Mȧ���*��۾���J�D	�?5�i�CE7�+��\�i�<�3»E��a�v��G���ll��Y7ۦ%�/t`��x]G�|���LHc��"7��ml�R��n�R�-��M��|����=fH�l2j�E: `ӹ����H۰Cj�F���ɱ��[���������M�H�j��~��+�Nm������L�;���D8Ǯy���������=�FF����P��c�[
$��1�ǜ�g����С�o����=��ر�[|��ch���T���n�z�:� 4���o/�X� c�g�MX�Tț�=���1^b�iQȕ��!0���W�׽6���ە۬kK�Ī �nI?<��U�ᠮ$2Wk�)� �؀r���?����z��4BsKmi�s�����hJ�f��g��×�
$D3U	l�)��<a��owW�f[��� �bb~���\s9��>��%�V���L�~ڼy��.nz�>�D@���nT���ݡ��>j�:�OJQy3';��������P�����Si�A�����u�>2o���n��?�;P�T�
q!!&��QS챇�*��\�����>B@MY�mE�e Ɩ���+�B�A�['�/�+C��~��B���xR�"��RA�_[�CpLd��eP}�];��>]��ۆ�����2D�[yt��߇lpmte�9�B����N��%흏'�\�Oyn~�K�c#'����y䁴��z-�Y\��0Vp9�<��Gp��Z-i�W=fE�����;'(�4�z����+�
|����P�W��A�}�1���y�L!_��(�ՑmVJ�lA�1�X��1q|�/Q�l��~��23��"��od���Q�FGv3|�p�)�z���2����Hҵ��Z.�/�P��$�e��)s�+�D#ּ޴�r�m���*�GU��j��ٽ3�t����$؇a�p�����⒭���k��3��P�ƻ\VD��S��aLXaEA�؟D�]�0Ϥ|(���W�.�b�����t�m����s��<���V[}��e�c�}G�6��׫���t�m�����Q/��#�H�C&$�� ,�8G�Y�EސdUA�_�'�z�v}  >� D�S[�|��R�l��X*d��_�4g$^5`��Zre�C��o8[.�rYׯ��|�譎��Z�:�I�2��)�ʕFy� q-R��f����i�(�orE)�1`�����1�ߞYl*}����Ox��3�$�&�U�5�sP���8��$�W�.@
�M�=���)���0�k�kb�Z#��f�2��s���ސU&ô��$Y�?SA�����(�2�Y����V��c���I���M):�a�����'��6���z7�AT@���t�x�����ײ���!�ἅ�ՐK��M���
[��,�7�)~�	BX�	$���+S�%~����o[*���� ࡆ��o����{��h7���	��ks�`��nc*��hf��v6%Z�Ruq��z��vd�C�ͅ�U�����.��#�\�?�A#l�|�/]��v,N?�]���")�x�@UoY���c���O�F:r(px�Ml��j������3MD�V8���f�9
���@	������xQP�@�$�_uRو
Y���h��v���E�G�U��[��5g�,�᮵��d�R���b�fڴf�\�'f�֬���kǖ:�ːD�b[LV�GO�i�����/����f�-�0&2�e$�s�����N��'�L^G�Ӣ ��jd��uhsakAk�C�����
�,4)����h���J�>��ބm;A�C�f��o���#�H��q�R�˵73��x{��k����[�֜)ae���|�cg��̝�r�-�-sN��I�S '�١w�k���O��4^36�檠� ��Zk7��f������7Q�&#�}Jg?�ny���@��}��b�?Ǭ|E�L�|�M�<E�+�.o���;z>��k�g`�w��۾
xR���_v��by�\����zg2���r��G'�(��2�QY���+w�"���H\}a3�=��YO��g���/_z뭊��,97�1t(�<J��f�i���y� ��pNkahA��)R���e����rL	� ����0*�`3�x�܏��=Mo�
ת�N{V�.��W�֪(��L�M�9�"	��n��Fs��IR���?|�X�8e�i���O��F/?%��&ldB�z�/F��I�2�Pfn��i��ߊ`�6�lz_�ʜ�>D���؊֭S��L��-.yf�y�vվ�����[�v��\6R�~I��{��U��8o�,Peބ���n������̅ͽ؅c���bK!��1�Gp�OR�k�aҒ�|��8����ȍ���9�7��/��"��Z��W�N3��yf���I)~-r�1ԣ���� ����Ǝ:L8:=0�x�*9~4�����J�V����P&׋�K\Z?⣬0�+(Ǔ���`ݲ�ì��S�	���_]�q�ff�+ �7��,�X``-&GM����k;g+���H5Ev�w0W��E;/X��4�cV+B���'��ho �m:�|i&x�Q���v�{�hr>��)�/MG�Mc,���CV�	��/!�OwNdƢGV�w�b�N��fjB��HO'����t~�/J�aY	";��"�!��)�\t��Q4����v'1��M�������EE��yN��>�CV��:Y��q'�k|b�#�#��g~qe3k��
���I�$���^�[���'��TVjGn>G�&̭���;��� b6�O�	����4��x�$'����-�Y1�o���m!��F�5E|/�d�.��+� ȘdAAؓBT+�;c�l�52Ȥa�����D��?�?7�4�b��`���Fo`6ʴj��=Nt�ˮ���zi�`��H-�FFXVM�.(U�%8�Pq�6,�,�U#��a.[��2N�vS�Q�c�r���I��R��g |�~q�K �� ��O�G��en��d8Y�&O?�[ H�
`瞴d��f��⧃pc
Q�͗�'��Q��R,�H�|7jZb���#�Xx�ZM������P3�W)�N8����أ���z�X�3����s{��`�ή���꯽���B���G�^�pNJmg�g�M���s�B���o8#���pi����(oy��H�L��$�=�d�A��/]/$�N��7)p�<9J}�>y�C⊏81o?�5Q���4♫������'M׼+��@�OS}F5`n2aG|�5wėCL�Ѿ�_R����gW0+�y�'黎���^�7e��S�A�"� �E���Jw�z�~��9��(zj����y���F�19y>]��o#M�3�t�wzy��p-���J*?}<���H�3*.�H�Cn���U���,�D��Dv�l2��ĕ�	7sY�Wm��!K�m�#7+i���
���}0�������j��6ک��X��tށ�:Т�Al�����,����������5�����?"&��r8�Ԍ<�Z�%�/�O�����+����������KT9�Gl#5�e�׸�$@,���K�X������t�pC�\se[@���4���U������A�����;ܛJVe��Y��04��L�ݳ�JR���я5��Z[.�i���A���2�id��q���?_�O.���r7E�������Џ�
�Z����R������p�U���}���䉣�)�r(�`6�Gd��؁N����2R�sY���m�0�(����
��/r�bP�#~�o�B�/Q��"�`#N�w����b�Zk9"�����ZAI�&~AJ�������.7\�a��S'��|�*�%\T�$!����Ro�q�q��n��vM���mQ�e}���Gv��>�Aƍ�q0���*����Ћ��F�YR���;���K���m-���H���DI#����F�?�T�������B����0�FL<�52]�W),z�Ո~��Ck+(sY��%z��P�F�Ԁ�8F%EО3�v�]�/g�Q��O��5a��p��ϙV��ml8$X��*w��L�k�6z1�9�����v�S'4.d.P`�T��e��T��?ah5��r�D8ex���o��B$���
���Սv���۝^�][��������o.�+ǔN�ci�����ղ�L@�h�Q��d��-5�:����ȠU��^
zڼhUUr�><�����.s�m,��V��T�J�d�}4u��%K��y5x<���;��)|c_�y��S�� CZ�)1t��Bl�<C�1k��](�&����V�Z2W9Lc׌�t(|�!��y��������%��<a W��\�ې�~��K��9s��S�s͎�Q�_��t�u�m�96���5��JEd�N\7�(�� Z�w\���FkwZ������(�<�D�./]55𤳜�
�؉W[���kD�2����sx͝��E0i�83��gx�f�h'��	u[��U�)�ۏ���<^}�����#��$��,��=�J��gԡ��6E�3�{��T�;��4��b+>sI�V
�n�K�</�SmSz-�LB
�WE}V���OD�.���$vJ�J�Y��?��B�Ԁ'�(�uBf@�f}�G'h�`�R�u:��:e�%3h@�
\M��-���m� ��g��To����9_��������_�D��w���y���7'D����~�v@;�@;d���w�%w�����!�������6ڹ�0�KhQZ�'�����?�"7�b`s��������{Q�(�]�}UU՝�H-g
����`�llu��&k��3�O�RJJ�9v�����{�*���'���N��f�sS��5�VK�~��݄
�2�o�H�p[���j��˲|�V����^p�	�&찅_�4�s_^a��{b{ I^ڜ�u�4���֋Y�ߘ4:� ��Q�У����V��Ctr%�5Z�a.�2�ø�/ 1z	z����2�5o�n}����҇���Q^g��E��3��+��D�n]��Ф�'?_S�bE\ 3���{��,6�ǵi6��=swA�X�x��e�GL�q����:�ߨ�_��}��`u���Ľ��8ZH�>+��1z4��N�T��d`�*�"��3#52v��A���GGr�w�$�nlʵB�e���_�ECM��7��s,�v��@c[/����tM��$�D:H%b��洞[n@�_,e��`��Q�c[�w�Jg.�^o$���2�����f�ƺmb�+@�'��b��r�~#����h��2����iؒ�0���F73<gLca(CuW�XG� �ɲ��➀!4i9QO��#d��˄LϢ����\�ɂ�I���3z��u��]�kKJf���Oi���@wϹc�XP��M��gf��n�Q�zl��0��g35�UJ>t��,ɍ������)�����`R���P5��@i���&ǥZ���6��UɊ/]Ƕ#gb��?��>��"�>]��F�;��Q����h>
�4��D�sl��:�_}Wq�J�I�);�acW��Υ�m��d1���%ٔ	�*R��%��(A����>�Plt
d�SC��9��6TE8�~��A����<�N�װԎ����?$��)R�`ѣk%�G�D������V$$4�n ����4�@��U @��x�o�4�W��e��nZ�S��S����d̙ �#\�
-p=�|r����~���iA�
�����#�0��8AX��NӾ��X�$���6h�O몀*o��G#aj�F��Hp�&��jHN����T=�&W{,2�m�����S��4��I[���6p����YbI`��+3Q���b����}r���z��!4�&�J�D�ar��f��F|ȴ�Uv�H�d0�S�������I�,�Y�X�(�*�x1��:܁>����"�����L)S�C.��ξ�:��v�����G�����lL�˙�a-FC1�W��^w�.�'wd�/w9�1ŵ���j6cл�zVD�4kT�܁���%0��W�OG���cohh�7$i��0V"�I
}u~���On�����1��J�^x���%��Et -�R$R!�h��d��2eB��'D�)Q��O!��Nh���yIˁ(Nn8�W]=@�.���٬���o������%ΔP��5�0Y��-G$֏�s�;�i�޽v[�#&�p�AH1ib�h�H˃�����c�LQџ�l�;T�(Q?0h*MX���M������8:6���쳼��;���pE�%�W�����? ���#uN\�C����$�pɏү��͞�m��]�@pч�����>�W���StT�PIu #^����T{��?�g"G!�0�G>��+�Uf��201��E5�P��ˈ7إ��V�ir�eI�~ݶ�Qf~]�#���c��2x*R���d��o7*���Vߦ ���.�%y��<��j�#�b<��u���%��,�V��ɖ������l �8ql1,�u_�v��4�ف%��n�m�/'vGD��"�J��E5�F��!�K�z�R����k�px�7�`G˴�-�;����G��<�fN�D��k[ߋE����������l}�(���[')~C�����g���8G%
0���uUZ��@��W��3�WA`D���d��/5*��+/7Q�"��DU�1X���t��sy�Ə *�? ������g�6��a���Z�y��D}녜&�"��6����D|���I`�X�J��^��9*~e��I\��+�n�\�4O]X��"J2�|��h҇r\w�����t����Y�H�h��߷Q��+{�H�� ��~E����*V��&�lLr@�F�|Ul��+�
�Y�Ak����׸��Ŀ0~��q9�˥1�͙բ�3u���&N�
�Q �����ȳ��zvv�����K���o�=9h}P��9�4�4	���q�y�N������$�ˎ��'�#ֈ��ޗ��,C8R9ԥGGi�_��;���(x�W?�E]4������Ӭ@N�&`ݝ�bMu��D�ܤC���������cW��_�k��ve��V�Y/Fi}{J!���h�ˈ����sw�c �0�/��T�m�iHི�M�uR^�t�q< 84�E�4��G��!�+�׊L��hJ��M�0��ļ+��[Z��`By�)h���(qϮ�cɽ���q�7�߭C�w-��YBߞ�4��ϸ�bw�=��{���v��u2��$�y�AO <�u)ȭPY���H ���w�s���`����4!�g19s���0�����3L�0Bt'�Ye���ܓ9�=�m�L��1H� �m��K��R\���2�l��8�����W��P���ȵ@��t���MwA>Y���UlL�{?�J�J��+]�\���/P�.y��B8)AAs�.p��v칯6��ߎ��:�k��ƍ$����AD>S����b����[�a�!G��g�JA��RkN�\�'�4��Y�� ��Lz�N���'����"|����p^a#&f:/���:�(���OR��`
"~�m�sՄ��1E$��T�|������z��S^shNh� �i�Ga���٣�T�������+6��T�D�f����iavk�>�e�`�Td����TA\�Cu�Z_�c~����eRR�'u�9�iSi;�w�+�Zy�t������;�zeU����\�#�
��D�!��
̥<Z�^�	�m�v�����]�Y�*����$w_�8��)j	p[�懇R��ǐ{!8�P�
�
����<u]��v���bBC�fU9��>]z.D����,!zzx�5��b�=:`S馸��넖 �����D�jN���?�!��`gv����kPQOKlYm%�M�%@-�/�ˑ� ]��Q��V�e���Ke&l8Z�B[��&LC��m���*�J�'��5-�H��6��B@�"3Ke���$�TAe=�bD�n��D�w��i�ey��������"k���{O�ג-$��EC؁VuIV��r�-�޴F�Ѳ_L�Z~Jnp=|oDGs�S�B�vR��}'GR��|�&��:���`��ퟒ�G%Mr�e�8Q��\<R�m�a�I�s,�*
�Ǝ!�.t&�~�aEA.��kXo뒛�tdL��~Ĥ%����hbw�l�_b���8���`k�B�`��6k��z���F��a�Yz~���
δ�/y���Y]�(3�^w/7����Ա��5��E�	-Oz�5��B��C��lZ�U�2�:��4S*�ˁ���G5�"hjY���xΦ��b�}2'=1W�<��P�!����!h~q��%�\��_�%s'�Tj�gxG�Y�S�F�q�dG��hG-.)*r�ƒ0ݩ�f��7�|�!��H������3�֒� Э��l�e���`�㜪�mU3���z����R=AQ��R�dkW�փa2��tY~������O^G3:����t��}!Y+os����OY*�E&��J:���ۼ�7l�L�1�Ο�yG�g� ����5Hw��N�l��	8{j��7_5��>HEc�.�£��
O��H���-�AЈz�,�?��r�(Z����;|��fR�H�*�u/R	��~H���6����gz躛���r/V���ʑY�ZX����S�$�yT�'4;��F�n3�<�6�-�G�G5gɹ)eE��i��� �,�݌�̻u�|6�7��]-�T�%���7���z2�V_j7��s�
 ���L���jK��j/��8c��mR��b�����RAte;Q��N%�oB�]��M�š�lmNcf[�ù�a��e�LL)�5�!1$m�QB�%��y,�P+�!��8����=φ=��5F7H��z��&Ba�����W��R�?A�w��%cv�X�7�:=�3)�p�q�+Cm�ЅK��b�+�pbꕣ&ZN��J]�r|OĚY��_p}����f}��/M>��)��}I_�~��΍�X2c��	���[���b�P	S0O��6�\Y��i�`��T���fR}q\���{�@kh��l��\Nmk��VH�p<eCl*��$���U�vw .��� ���cԡ�W �.D0�/Z�J�'��+����o��NUwyf�����Ril�{����[:�_�P[?+T� L 0�$O�ο��xiq�iE4:'Ӂj��KKP�����}Ί�P)���Lo� Y�T��K;�d��<ԕ&�z��,,LX]!�݆7G7���O�wa�f��6��TO	��̼�I&i�]���TU�+�[�%�][bN ��Ak64*���؛Y�[�)i�Ȍ�N!�P����݂��3Qϟ�8�<�������eiK����㴟��Y�aL��+��̂>,�d�4��ᢞ+㪷j��Q�����"X�8��mj��[��񷚤����@o&9:���e:�l��"Y�7@Xh6��'C�%ʎ�h�Po�u�jύ�Eq��WZb6��kp��^�@�0����ͻ�.,v<nk$�}p�;�d ��딈�*o�xk-�h}H��j}�\���{���E"���W�
��;�y{.g��KU�O�D6iE퀬Զ�E�k�h8/*�*ޤs��X�'R�q\�sT�̈́�	��X��~���b��q�ߵ�<���=i@�Q�m0OR��t&TY�l��>|��K�'V��hd�*7����_��((�����v-I����&�	=�(,��(l ��Ƨ�������؝�w)����<����ԋ���ÿj��Y��Ȭ�j��o\�Kx�٥_/�:��˸�*���+H����w�"4(u-a�{�̓��3|֏�tC�I2w��cR�r�7��Qr���{_�WM��0p[}��.��%��]�!�t�⫔���Fӱ�J"v2�aC10P���vO�k'D� Il<#kPa]J
I�ڭ��6��+Q����W�n�[Cs�E$������pEs���2'�ܨ��3� = }�G[�q�������Q�?���`j����J�X���
\`ȳ�Y|-�td�59�`~ʪi�,�Y}�}��K"�:�UL1�\��}��ss��ЅB��S\��}ue�Y���/0P��(	���9�{���N�g�4�3��j{C~GUY1	|+���� �<}XK>ĢN�'��-^~%�N�� ��O�u�����91��MP�n����Z�E�~l���.򅰲�v�̺]�1�������ե"��21�(�>A9���U2�~w���S����Tir
_�kP&a��Xy�d���f}H9C$w?�eD�IgW�4�8:���K�vH��M�W�)��Eus/L�AO��.zE=��s���3f�MP '�1�	J�r��}�O��q��!��2��`Q��(nBI�O5��r�Ύ���&��<�M���<<���)��mmi���׃O�m4[�ݛ��×o��mY�p���J����d��	�Z).Ԫq�dpDl��iDd9Q#*b���]���O���2�l��E���e��S��BQ�\�%��5ӄ�&)�w����)�Bs�E���3���:6	���(QqU�A���p?���"��p�c�<LL�����Y��`י�ۯ��!� ��;lQa⡹u�oS_7\�b%����djx��	M%������<��Ʌ'7U+��1L�OK�� �T;O�*�������oQ�T�k�]���`-�b��/�����f�f�"�� 5��~*HsIF���DA<���"Hc��۳b11����D-�� j�L[2�J�&����b��?�C��&2�.�樇�"�"8k�]�vC_��v�vzo����0r���9��<?�t��6HS�u62���ܬ���I�|�C�r\KJL�����@�/�e��`U�@+>n/��
N�R`�sq�����q$Q��}�~|���W��x2>�T��)�>u:/B���aKb���%�D��-�{G��t��5#���0�S�B:�R�̄��TA%�u+�����V��'p�A���*���#e����hJ����a�K�vɁ|o�`21����ACi&�8����q��qTTu��H�
���@����������UB����񖯼o]w��*nDA{JGU�_-���
�=:���a�Z�?m�Z���|�p-G�Z��T��?�9#�~m��(]��u��ʰ�A�N�1�I5�*d6�Sgd�Ll��+��HLe�x�Q��mqБv��2��s'TJau�C
v���w��b�
������is/^}�^Twz�"!,e`n
b�'�3�:AbkE�+�T�6�\0���U"���9����D��8�ۼXbT�6�cD\\6o�����_�@���i�o:;9f@�����#)RvJ�q<��Jd���G!g}s���Ύ�0c7�H�����LV�1\P�R�s��g<ݴ��L����.*(�,Aа|͖�b�&�Y����6�{���ލ�d��Ⰲȁ�� ~�Xf��Ue�=��o�� 9���6����u�7���N�;��Hf��D	5��'���Z&��u�m����(U��`�3P�2KMIc��k)��찄�;x������e;3L�QY�">
o�X� p-�~=2R�<�$E� ���lVY�ů�hN�'`��PL+�~]��>���`2i,,z�B�Ǭ�����>� H8Յy�1FG]!Ҵ��9�1��NN�S���$;uA�"e([�����
|�������Ue�KeV�)- �6�w���cA��L��T��6$����Ļ)�j,��D�`��\V�u�(|�!fŽҳ��R}~F�"c��d�B�#z �
,�/�(�"�u�1�]�����1F<�h_bv�-t�(č�R9��^߁���<��''��9�-�~H$��T@i��KѠ�}@�"iB���<��+�	b`�����}�9d*J�~\ e�{ѳe�I�W��^�QE�jF+�2��o��C=M�/��������+{t��ѮƣAֱ|Aw�����X���o"��."�C7e�(!�!���?�Lǜ��	�G[�c�tś��RRt��F��:��wC�Y�eX6�h+f����ൂ��-����EDI(Nk�����ѳ��0:�� {g3t�I �u�T�I�e��~-<�ܟy�~�y����R����tu����h.;��h#�5������ ��[ژG���:��D�0����������}܄e �1Q	&��?���PZ�����>7��ҫ
ȡ��jx�g���4b��b��&_g>��y�I�C�'��O%ÈZ�0��B��_%��Cҵ�1~E�����!P�I_�>�WSA�G��d��b��WU,�'Q��?dC�if�١K%,��a
}ttP_vM�� my�S��U'�U�4/������}=ڬ�{��B�C�̉����, ��mE�^a��f2����Th&9��vq�j��`S��qhuc��o"�{G4�T{�M`&e��v�����Wt
����Us���C��X��?f��+�T6�E)��h���¹�t�����ab&�\B�8E���	ji�/���oG� �IM	sX��!�w���5��r�F�W��*3Bn�`���}ܚuE)�@�<�� �!�[5��6L����Z̑���g�_��������DA��&��Q��� ���m��������f�MI2!�nۡ��F�Ew7WqO32� )�����"0`��sԼ���x���3k頠����ȓ����i�����<��G.��0F�s���f�oIݪJ�):���c��y�'O/Q��U|0~���a��E{��I:�D���j���Vpl"eD�	`I���:��c��r:��52Á4���k�{Af">e�;!�����u������a���O#r����	M��Z��O)��=���0�K��;6�!/���v�/�NI�/�ͶFVƨ�ƈ����Ȅl�d�:������O�	;�A�GU�P���h��
�՜�*+og4ٝ���L�f{=��9Z��b�����~f{��)Sf^g�Z	�%���+!v�
$�����F\�5����Hc�E�B�v5�w@�?�;�s	>@Hܸ�.j^��_�W�<]|��b��S
O$��TX�};�b	��HXq�l���Ra�9������^�8� V`���^q?�}����)HCV5XY�������R���$��:��b���so�9�l��)+
�^z'���a� J=^k�[��(����������K��j)�� ��a?Б>П\���a�ByV�d��}�7N�l9��25�J�O��RC�U��&���z[����A�jmj�j䃫 "Zz�I����C�c51%�c���OZ|*�jh�+��!P�i�.�~�!?I��Ә,�ߩw�]�Ba&��D�����U�W����[a��o��ӯ�h�:۽��@��#�n�c��Q�l�J`��LiB��~Ʈe�����nn)�]��O�$4��a�6��+ks�����ϧ�L�.�Z���`4��}VX����W����3�n`��r�v��~��cĒ؎��x%����޼����K��&���-t�����fDS
I����@?
�Ƀ�Jo�� ��֚{Q҆*o�`��	�����ɉw9�_�e�-�ny!���U�Ne5�Η-F��������	�-M_��p!��q�UÓ��W�Ҽ�ٙᡉ��Cm)�ڒ��1# mw��-�u��<��A܂�c!}��I����F���5�����΃gI\��&�ju ΀�x�Vمmx���cm�@�1��=�O�b�����;�XG���y�75�KrY�6:E�?��QPx��y����r.Y��_��
�4�	'"�-A��x�\v��Б�yz����9� ��Mf��B�j:$ی�jED,��,�S̏@�6����)�?ᕼH���ħZ���T��m���b����"o���[I��|�'_�.A�`��=�v|d���0Y`�L{�+�����Ó�'N:���ٯ1�cG�E;%�`2{
\�o��7���}t4]~ϢD��?�+K�!¦�=��y�3�.��<7$�<�j$�$$:W%��ơ��ݷ�f��Z-kȣ�	��K1�0�!y�lDM��C��	4=ǒ����u�.�6n�+�����r�kqL�D^��?:;��ez�}p� ����%�i��$7٤��[��(w+�k'�&���+�?Z�Jw��v*�.Yz�t-@�R�ӄ"���~c:�׋��RB�G-�@?H�35JXejbe���g.�ml5�a��<�Ι2�:��@a����.�<�`{��V��N��=��dcMzǐ��\��۬,R�͉/_A{�9�
Hj�����H;⳵!%�T��r>�g��#�DEW��1$i��EN�S?���W{�q��璚Hc����;ӲmXp!��xq�?;���b�㐰E9n��i��t�
���X& �,qQ��Q2�2���w�� �7��� ���]��SA]���_ҥg�$A�>0�/@X,�k�8�d*��@�h<V�L�F�#H��%�v��X����G�.�QW|������>rfE�V�Yb��/�.u�GM{���|��k Ԇ��$%��Qk��������Щ?/k��mj�u�2u���ŉ��R���)��e��LFxT���h����Ql;�9~�Go�	�Vطz���ƻM#6}>[q��EMc	������D�̵�"�z�}ǘ���v[�>nSHk�p�fݹEc�<I��2!�m����q�ɫS[(�aCC�{S�4ͅo?]��u.�G�v�kwP��<�H�/�������t����:
8��"K�3��V5���,�6�HM*RA)�D�u�����;�Pk�}ߥ΄��t����U��'�_��h�2*�% ~PZk�w��e������T�}��m�eZdOܞKV֣�O'b�<  ��;��=i��� _\�B 3Oe�w&���6�@��K[_�ꘚ([��,���XK�" �*<lLR��8��:|��u�( �y���з�]E�I�-6L򼪑��n���<�-�m�%��cc������h�$�e�ڲB��G?���U<h���o޽�Ơ>B�)�j�dC��v�˱�&3�2�sy(�|�M������ڎ�H�&;�!��~`�&}�z?���5��� �LQ�ǒ��63�H�Tv�Y�_ˋ��\���8*���TWa���#E���v�S���'��?}H����S��4�~&xB��i6�9�������\�s2N��H�hr�?^f=�x�U9,ϣ��������f��
��2��y��Qf-L�as�g�G�C�0!�f�y�!�-��Pd�}ï�w�T*]�l��B�;��=q��q���9�`��<5�\��玢��=�Qn9�G����a$�������e��?[��Jz��?�� %S+��,^��) +.IR��s�x���+_��K�	���b����UJX{��n���o�{��U��m7�Rz��M�	h+�*�C��<��d��^�^c�2��L�4������Ʉ9�|-�N(|jO��@gڿ�zD��"*_xۨ� �ɩ,�J#�UqU j:��m3
g���V���g�f���bT��u.^���
��,:۪f�M�8�+?J���y�-��,�D����zA	��>p�}U���(���{��	����?N��4��r�~F}�]��yˁ�8h�j՟���Ӿ��cq��D�������-�w'P�߰����N\}������1�S�R�X�j= �Ǽ��k�S}+�Lʳ�k}�o̳IU���"�0�܋N��������ͨvc��!n���N�>�ou8�o����8{a�Bd9�O��a�N��q6���s7wX�U�H�)�&������[�{��%'��2I{-6J�働"o_��,e
oN�O�+p8����`�CN��2��܁�P�l!�<A��o�S��ZP㒾��z��8c����?�pG8��fbCl�J��v���4zS'��U���w8��%b�m��|��j�Jl�M)?��Y�SmI  ��Ԟ�'�b^n}
8h��<1s�60^F	R�҇���[��v��L�.��ZQcty�xN8hp���U�<R���g%�[Q�k݈������܂����o��� ��qkfnq���=���)�y��V"<�1N'��oCs�Z�Ŧ���up-��f�,I�R�s�ͯ�?2~T|Q$�$(�oxG��L�\�?�A�ɳ��a�뾞�|"����,���=o��]g��#H��<�:)�����CE�T�V|��$�]�E6����k��tuFt�����D�Y�"eG�A$���@�Dx1��z˙%	��~d���گо��ϐ]���N�qM]����8L̔H� �k�� ��Uʹ�g6��Vڙ�e��9	����U��l�ȏP����P�Q��GP��Q����Ck����'+�͔�Hm4��/G�_z�lm`>H�	ފ��kG�~��"+�UCc��8�y�LÝ��Ϳݯ�b�4��{�o�9���1;�='�j���g&`*�	��W���	�؇	��UWE��c��ý�@�8ڤ�w/M��?���sM�K�6��Ī�e��H��5��L��{(L8�����&�{|��~N<�y�!2��c�9��~�5�󲡜�J�]Np^k��ӥ���$t������N_|���X�G��d��d���u}���r��l#�Mbш�ź���D��3�wE�[��0�T���� ���ۅ0@Ne��	��%+��诔:b9��0	�3z߿d��tfm����$|͊��u��1m��~��gVl��9���'�X�Nj����u`3������;s:~ۼ����z1!9&�x��� ��S��|��Ix�����6Vw���9��cΏ����cҐ�*���5w�O�~���j��D(�ҹ�܅���/n���/�a�pqK0�|�s�?�0��/��"&�0��<|��O�pc1��M�V��L}��bfW���Q�7�����7ȅu�R�OY�����E�i	P�����t����綠� ��_`ٛ�y��Fi�Eb�g��׸C�e+��-�,Bm���V��e�b��?vYV3%�J��m�6��T)'_i�?T5�_k식HAO ��6����$T�]�����ǽ�V�	�#��E4O$��x���egJtB�aw��F��u��B���r$�E��;*z������:�~`׳�Q�Q���f�[BF�\�B��[��<-��~�(n�B�Q��񁀍QP��1w����y�:lk� <�+��JO���k8����A��jJl[�}ֲxԇq/���z�n��3��^�c�Ɂ-0�1��ܿ~���=�n�P��t��se���ϐ�7=���%ǀ�K�Ļ����^Nr.t�Y��K�md���3�T:�v�Xd-�����lu\nޅo|�TF�d���l5�X��4����c���j�l!��'r�C���×��\8�A�\��	O�RQ^��&�u=��8"��5�s���'`
�!�RS�ލ01V��L��[��7�5I��5���Ju�&�ԄM��L=jq�E�m��UB`�M=�0*���AL�R�NgJ�(Y��{b{��T�(��˓8hA��i���U�����F���{��|�q���(���dOg�_�sEҌ:ڰ�6�}IX8І�!ӯɾ�����Ob*0�Φ�}W*ŭ�84���;����.0,�u�Tl�p=c�wy=d�����Im(՜�`n��#�u��cގPrr|�?<"
99/b�uHC�sn�(��4+v��2S��'�'�8��"ڮ��&o��/�4�Q��粂~��C�O\MH�e)�>�:���Kf���"�h�MH�'��j7��ͩ��n��3��j��8�*8A���T`���k�|��;����@���%$�]Ur1w�0@��NA1�3IU j����0�M�z�{��S�l��	�6u�4�J\r���)�.����*�Ø�чz�'�r�zg���?I@��Ay.j愿*qgO`�rB�df�5t��t��u36����Nj��3��P�(���=��Z%ue�H�:g�j�\�__���RK�\v��/в���uZ~$o�2��3���o
,�^�����x0m։�2�z�Ÿ/[��%��[�����(ԅ��@6$u��#g=b�{��Y�2�$�8>���g!Y���۹շ���(���H�
�Y����~���P�F�)��`w�ؕ
Y�����V8�)&gE8�v߀�I��O�@2'%�i��1$3��.j�Fw�hZ�@���d�t�{1�=I������Q��y9w7�f~Z�Ҷ�_�2��<��"3o��h	hsLO�N�rv��pԉFɋ�$,p�{Y�QH<g��qa�=�^_cE�X�?�'K�7%n�и�c�D��$�`D�p&%�'��#�Fl�%�gx�u"�!4B�%��)w��m>�.6y�X60<�V:��v1��vB1-w�`nU�o�����~�ُ���?j�]U��!�r�ɔK'i��#�Z���۷Ca����&�,�����͌��4&�sf8Ax����K���WA��,���_cƲ�߳�5��D���ۗރ�|���fZIxEJ6�ђ�'b���`�b�6��+�_ԓ��p����cР�2K�G����[R�6�W	eGq�\�{.9�IA�)�N��<�tx5���}��~k#�J@��T�_���Q�����7��gu��8�O-�  R��L��@�6k�Q~%^=�Kւ��k��r������=.�͡�%�HCW�'?}D�؎�8�`6��`������8&�+�i��%o�]���1�������b<rpް*-V����Xd�=+;$]�9P��ܞ�"��fHͽ�i'�{'J�V��Bx/���i7�z�����Q��dt= ����f"��P��Ό��ڑ��)4��kd�%���(����u5$��#A�����[2ܪa��ӣ}b�W������)�q�a��"���Gƻ��aǿ5�Z�Y�FA�0��.v�"�Ou�,K��7yG1��}��vғ��ΕN�P�-��yT�{$�L@�sA��DU:Sַ�B��).1Õ3�MJ<�}:Bd]�~d��L'�"Ӿn�Fp,�$B/4���m�7s�2HߑV4�������}іqY�|�q
.��܆zn�#8(�8l����6Ҥ���F�y@r���J�G��l���r���[N�E����;�-W��=Noѱ�8�S^�|�
$��������SU�=j�/p� �D�+9�o�WB#y�e��Ys/��W%v���\s�S��D%�|��y�C~�Y��%������iˋ�K6Ұ�K=hO�~��N��l�K�s�*�����|��܈^�(�����c��w���'�A��3�����"��EQ�3�FN�	���G���UU�����#�n�g!?�QE��*�)�<ԟ;�o��������E�ܫ��nS��������v!��T�dW�w�m�L�K����I��sa�?0o�E�d��H��~&��*��#��<<ɋ�w�=��~��
 ^�röZL��g4�k~������m����7][8!te�YOi߾�$���Q=��Ly3���֌�G�F��5CV�Ti(���h���8�4��3)�Lk��yj'�� ?����C�>�����I ��3us"x[�ot\�1�ub�(�H������>rb��Z��Pֺ�&`؇ Xɟ�3�y��1�~���H�Gf4n=����Koׇ���o�ʭ�V�~W�236^�O�B������%��(r��;��s��s�\�Ыz�?���h"���~�9B���qE_�u�d���`��	0�1�e��H�-�(�'�C6�L�q���}##��\j����a�תcjf�ǿg0*����у�T�F�yY���A��`Ф>	 r���Ch˺�;@�1�vh��!tQ�"r�o���C�s���C{��������L>�c�C��4�Mr�2�0�y��u�9�OD�dwj�C��V҆�e!
���[WH-oۥ�A��L��e�s��
��ϊ����c��BؽC�?	��:{J�'X��R[s?�F�hC��Vƹ�n�~�qk�A�����=���W% �G�/Y�cO�lbkt���Fj��MO�ea�i��jGX2G�2LD�5n���ne;��֦��R6����8kl�
P���<�!n~����/-�K�nw�bd����H:sx=.Z֞��NK:֙/%u
�sdT>(~��ǣ�a�
�z����%����Q�/H��S���8���V����< D	ڳ����F�2���ꀢ7�"}�H�+䶫�A˿��ֶ���i����1*�w��r����|k����b���ړc΅�PnJ�O���P�7	R~#0>Ç�a�\�����}[�?��m��v��m���K�X��N1�[��9���ޗ�@B͍ g�`t�sT3��'��-�,�xbk%ċxn�}Fb����:n�-p]eȎx{�L�7�]��u�����6� ȝ����|ºo���n��*^���� �0t�x�y.��R�a�OqH�?���Q����"]���@^栙Ή�Oq�jP��n ���P�'����Ef	cj�U��Z�ep��/�[�M���kC㩉$�n��w��/��3���{Of|YQ��,S�ҋ��ʥJX�Z*�l��*m;t�.(U9�}��� �h�;k��dyK������KK�[a���!��K6�1��]g��+���65Ⱦ�Я&�n��|�@#�Dٱɳ��S2�]��m�������;�qt-r��J� ��)2��v��+�J�~�I�o]>�!�X��u�E8a��`���z�l���M)\��*�:���y׎>��c��ˈC08��w�C�	f\��aǙ�R�q�G�l�^`?|!����pkz�&���r��&�k�[e!q#�yqߥ�8�͚S��@t��G	�b7|Uwz��� *�O(��J�Q$�}U2��>���DqkT!�
	ߏ�?�A�*��t��7�"��.5�txqHQ]z;��������@�`K���1��Ƃ���ҀM��+lMz"��iB �c��ϑnq�&V����`8(0s|��<�)��gW����;y���'�k�=���mh�E�T���%�NP�B�u����c�PeRK7���^���L���FϤ�"R�X���&����Bt��w�<iqMɧr�5b�tv�=�U�P�l(����!���}�����$�w��D�J�PJ�a�]|�M4-��wu�Vú�p�JE(���̴7�|��@�`�L���@M�����L�J� vDם3�s��w��>��$0�<\�IqR���P�-���d&j2�ŀ��>�I��z��4�GH�H2!�Iez�,0��(���n�<�L�0>�����E��V\5=�YVn�����mQI<2�燶�+O���P>�Z��j4	r��_U^�M��^I�G�1[��v�u¬�N"b�����o�L)��\|�������3���c(Ϣ ��ڃ���}���E�((˗x���ly�{͸<�>���t��C����i�S� Ћ�������n��0�J��{�3�c Il@�o�lp���C�k���8�ۮ�:�@��m`�c[�9k7B��NE�Ð����,uW�KyӍq����Ć���{r�,GϽ�[�_䣇�M��3�j�|�1�iy��7�
����� �i_t�	�{T�;xe��|��~�_�L`���R�:���j$X���X�;l!,]Y"璨��h"rn�jwBW����.����8�qK��rc�_O�9��P��?.]������{u�l��W�=S�v�	��jG��"M`3؏�/�:o��)�;E2<.����l�͋Y�vbN�$j�灴4i���8�{ ��|3�>I��2�������D�=2h��>Xt��ݻ��Ȉ��3�k�G*�=�p`[��WY���{���T�@�ZA�-D�<�@���_��VBp�d����pF��YR_���3��tίt�)_nY�s".6f�jj+u ?���b���p%�Z�c��9�zڗ�z��N)�a��-�b�@g������[��sx��qRz�m@�R.�ݲk-u��MSj7՚�$��k�pv
�M�?P��4�N�{r(���<�m�\�el�Xl�k���#A����|�&|�x{^�!�k�嘐��:].Y����A*�8߹�53��l��~�P�_�R&12f�Gȱ3��|@Y�ә�~k��!h0������c�ߵ�~�ܢk�P��%
����d9_�p�P�L��*��^����m�mJն��v���,�A!
�Q
+��H/gPdA�<}��#��6��V;.S�_��I�P<����obfF3�[(G��q�f��GK�������Y�����MA�J��l�p,�L�J^q?JVi�_�-Fx.�E}��e($²�/3�`�կ�f§,���#&ؼ�r�%�m
nX��$ѣ��3�ʧU?�ÎE��1�=/ҙ�������ǧ{q��M�,Q_K]�p0[ާ�:�_g_l�<�hIӠs�F���r��u��Ϊ�͆��(Vz�V���t�,Oђ���Ҩ�8˝����������+h�6�aE���X���.�Y� EN��]װ9bD8B<���X�!�%J�dɍ�3 <�j�"O_�+�PG�Ʌ���aFŷr1w^U�-�4�U��2�h(�xmwY (ݢ2���L���2����l����ۘM[��L�ƷR���
�� 旼�\��|��ݫ�e���$InJ#��J#$�Oם�U5м�Af��q��� ��>�)��ш�o[�^�o�:[.��˛tJ<a]�7��iƠUQ��+��v�I/��z-?�"�
m
_��$=OF�L��/{%�r��D���w�Uz�I�Oq�4���Y�����X����	Ȝ��g��5����4�^Y�'�$��wsSc�5|[܆��7��V	9��v����^���iFD~9��z{���d\$?�NԬ�|U:��=�S�q��҃��\0��N|!ֱ�a����~�f���ZkC���'�ܿ� ��?o�a��.@D����B��h��(d�pAۡ[��j�zgP��K�}��{O���s�����/Us<������T�l�D�H���u|�ϯ�1��>'���J=�?���Ts;�y�䬫�'�3ee��j+j!&�꫚��pƭx?��|��@ *���G��s��.k�x���Kkdx]�؄� ��\6�G�������򭴐��j��H���e\R�X�R��2��l��2Gr�҄G�J�7n;��1.{�,9?$��{�qD!Lp�u���QXH��H��JF<��r ���On�RX����5�B_	UnW	dG8��j�DH���nd.�^��_[dln1o����I[Q�W�>�y��]����:�]9��ڏ�A^�C~[��&�����y\j&�#�a�[��m1zBL �zl�����ߡ��ܗ���-qr���u<�ڝ�w�}b;r�Z���l��oG����cK{�⤩\���z�i�/��^5{C�Y�����z�sT|��6���Kܟ���>�����v���ykW9����]&+x> ��7 �m1�ڡ䶣����쐩7[��Lͷr\��2��u���}K�5���E�4=��.��va�B0ƋԾI��C�a��
=m�-��,�'��~gI��Eڎ���B^0�����ϳUnM�	�����x�NJe�^Qb�
W-��<��u_��ጄ@�J��5Ss�&�a[�OR�R�$���o4?{��p���އ�e[{�A�%ٕ(p�Sl�v�Q�Oխ|29s5�����ũ(L9(���Q�W�
f}��A���I!d�25�bO�c+3������8g(�S�ރ��9�\{����=��K��Q�c�>�T��]u�����	SQ�:�,gRf�9g^�+0���iNi(=�'1��*��%:?dF�8��t�0M�:����妊
x�����'+��2�;q�����<�Z�93�Wɝڂ���š�����,�H�9����9HT#>���K�ݹi�A-Шk�%�u�|��'�5T.]@a4�����x�M ��S���U?��Z�4�g����U��mڥ��l�o���2�ZI�\�X??�[e^t��:�*�C�s��?0A_ �"t�H�z�$��e
\	!��ϼ��r�MO�5�)}Գ,�sѠ��?��	�³��0��ԥj��4n�Ý��l����)��s\t&J�L�4C�߇�	�n�z.��1�J��}��^�d����M�_��g����N�&{���j���"�n4+	8������.�i8�wR�o�}"�؉����-@Њ�W�����VM����gse�o�Kt5�h��\�Q��glˊ��˨0�7`pb�nƐߣ���������wO��U�v4H��:��i>��u��S`�	X�m;�5V�û2�v���r����A�`p�6Y5}���E�}o�I�Hak��T�dX�WPs�h�l���;�h��W�Mȹ�s��k2X/�P�����[�q ���mhOэ>}����p�B��[p�x�@���O��b���~,d�t�ǶSC���&���gh��$bfb���c�s�w���c_*��?�NV+.�;u6>R:�ePn/zh�� ����}Z5�%@X���lt"bZx�<��҆�d�R"�Zu��)42�I�Mw�rW�=�]U�<�2N�7����RP�*���e���`	�k�m��+ܛ-���>��*�0@�Gb�U�N�H7����8�?L�5��ۺi��o��Բ����ک���v�e}
Ì���X}G�%gy��j���7��;�:X�1^|��TX=�q����K�tm�������N���=ho�qld>>sR��l?xO��me�$x�������&���T���ELz]���A&^�m��WHo�ũ�ɟ�����8L�3-5���7t����$8�J�ת�����N_Y �a��$�B�#�)�7�.U����������@�^L�*���ER{!�4_��(�	3M$9!yIqoƑa����q���Cl�8�P���7��1��P;U=�bd0��a�Z���#�[M���t��)��{�	���=�����Y�����b�� U��C��.������-&؄�c��Ư�ey���͈<��J D6����ˈr�ߟ�g-m�'{��Q�Fg ��:�$�]���y��@�3�����Ex»�$�i.�	p�L��r�pV~��(�����j�N�@5��J.��<�'|Z����ӌ# vR3�G-�[ɚ�=y,�'Y�5FB���꒏���т�j�/�̓���3(2�LzU]ߵ�T�~/����|gG��zB�rѸ�?F�~]��*�+�HTJ7ER$̥�a�e�t��S��j�䗋*��;��^Ph�f�V����д����}�>����vJ� Ǌ�̊,�7��ܐ9/���o��8�{�d�ҶQ�	)�bt��9�,� �;w�Gg	�O�î��
��pP��@�e�;C;�t"���PZ	N�#��m��YE���{̜[����?�&�8~�خU�(�E;��I����|��*��9��_~���8b���E�
�Q *�qX_R�`Hd�Lx�v>I��,j-ǰV�=c�;'4:�ܽ̐�Ug�[JO�S<;.��A�o��b��֗z��/.��<��rq̙-�X��<*�͵��X�L������;����CvoQj/�7�vysv�t���8����Eg�ǿa>3�v:�s�{C���u��
ώP@��)loq�I}�.$�ܞÔ����9v%����S��t�h72�f>U�%��g�p������j9�l������+�_N�n�c�#b��� ����]˦k�%gs����{�d�.�l>��uزg�#;�QLr��)g�$�\�o�k|0W��V�V�N���öхb��t�w�QCS|���^�Jk�6����sb�����:��U_�����&��&�(qt��F_g��m����'Ϫ`}��'k	����VS;�$���&�q�\S��gZI5-P⪺DD����� �`�-&�ɡ5J�G�5&a���Z�Ji���eTPB���< ��b��	h0���/!�]�Ac��0��)sr���,a�9��U�`ϊ]=q���q+��<U�L�8@L�%f����KGq�TM�c��<�z:r�bj�y�_j�9������=͵"�=�0o���R)�L�:���#�k꾋�VV��X?D�٨{F����Ҿ���:& �@Ω�b�0�L�r?<�lZʳ�Ub�n��W��G�� �kbj� �@_}��"r&��`j�F)�y�W6T���D^�~��࿥{���{�pս�|8�ʃe������ 0���d�^�.��z"at�'�UXڊ�L�ctb�J�B:O��#D\)�0�����M�2�\�ψΒ������v�Iis7M��15 n e��\�D�~��>�w�}8��Ƀ�X捛�)	�D�e����f�g]�C�R#%�sY/�D�ʁः1f�� �aX��~2�����q�v �Y��D�sp�|����y�`��1ա���j���V����N���i�[�)������K�m����(�-�����ݾIfpʐ��v��3]�d?�ˑ;"�)A��	Zë��&�Fn