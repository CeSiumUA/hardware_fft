��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c���bǳW�}N��g:��-�~9�R]�K���&6��q�
�d�d��a*���}�GPk"��uA����u��NzII�9�$�%��Ҿ��e���J�_��){I���Ґ����m�S@<�����v!�b��hA�]���L��/�P�e?Y��Mج �]Xٝl�V~�32h
,#p%�����ŝ ���ꜗ>����Va7J�@���M��&�y��#���?|;?�#Z��!�Dy!B7P���\�� RK7�����mZHQ�.�U����6y .'����}#��#���{���
-�2��+�-S{�Q@Y;"�w�g��Dgx<���m���J$2_[�C@���/���%T�qF\F��G���1zK8��1Қ�-����Gy����(�c��A ���EʚS-�~��{�c_}�3���r�G�D3J�J���@1_a�ê3��y��E�u�I�ZJ�?�SJ���q��Z���b}F�3|��t"�f�]�R�9N{�Z�N��I�BYA��
~��կ5�u>�*ԁ�E�#�ADo*cb��s+���l���N�(���sWjZ�h>W��|��ƻXYHf�����[�tՄ�Dc�7���1�3�ߜ����nJ<�I1�����I��\A�3yhY�A���h��e���P�Dh���1>���c@�C=R��#��E� ���#9[$���l��c����_/5�ݠa�o[�9Q�իF5���h7���yW�KJ��:ǂ@��%��a��$��w��;sz�Y4p>T��ź�oC�S���tM��ϩ(D���Ø��2���
�V�Q���ډI۹w��Jť�T���0z�`t���5�����؊�i�����i�Ol7�7��ު��y�
�=M����A�\q����GJ��v3^�R*p~6�]D��V����;����L�ڐQ����tH�3�F{����"P�Lz2���@C��*/��u����=u�m��R�vW�����D�Ƒ�d,6 eMn,f>�����C2y�%����k}��р��Ώ��r�A~���R��s=.��ykf�2�'�>3�36�0��a��[����5�A�>��A0�`��x8�*�#����[�8���w��phY��P�� �ޫ�{�� m
�KR�d�S�0���ƮU(	3ߵG ��JOC� i��Pe�����"@?%�����p�ߕ�^C�JB�t���i�{Õ,�;�Q��6�bؘ��`�h3 b��l&OE�K����˃(��JU���P_��2���NJ�>��Tg.�=s?#���[;��=��g�/G��v+��t�ɿ<�V؄_R�-Tz��ԍ���aH!d��kL0 �EFb~�24d �OKW�&KaG�t�����W܋�y4ac%�ol��{7?�Z��<��`�E��S��r��ϔG���b��l������Bz	әV�ZY�9,dK/�us�]��9�_(o|���q���u�y�V�ʜ�*�f�h��*~v2�{K��;'������w���"�C��6�8Ϣ�K�+)�sR|*;��i4�h�pF�9����� �<~\A�7H둃CTG��Z���O�n���csA,��������Y��NK����I�#���:�S�)Z��pxO�����[��׀�ϊ�d�.��al �����0�N.����RU�����iX�[g��\���QE�H1�0ϑ����k2i��4,����`v�0zI�Ł\,j9^P��K�w������nF#���Fp�U��f��M:�9N�(BR��Fq�Sh6!p#8LE������%y�D����H'Z䮆vy&��?��̑Jt�=��ݢ� �hOo#���D�,�w�l'G=3���#߻�"�@-rN�7���]uBA�H���c�����#��� j:��:���Q�'��C�"�'����d�ڠ�Ϫs�}��h�Q��3=�рfI��zb�$WH�
q� �j�&"���1�8��㈽ܵ5):��7/m��F��&�����@'������rE��	�"���O��R�"�Ɔ����P�� ���T��4b��dL	����1�1���ʐP�3�P�'��W�GS�'���:�g��6'�K��7ֳc�7��k�{'a͐Ҝ�!���.�Ka ����N�~�\ ێϧ}��)����xw��H�E,�zg���N�^����_<�Կ�5�qf��{�5	�d�L���l����2q�mG;�Qm�6xL�'r�tT�0s��(�㲟�(��<E�qzrC�y᮹6��Чߒ���yir?��I���-%ND��Jb8�rSS����/m���pв�)�9j\ǽ���Z��Q�6�
�����#sն�2S�~̸�}aG��.0����l�z�Me	����P�T�Ͻ�T��I�;�*D2&�4�����<���ގ�0�	�A[O+'��-��ݒ�z�����[��/���2�Q��]b��K���r��oͦԔ��6���F�G5���������]��츃8�{�����wRl��0}a��]��5oE3ޜ���/�_�#����f��=L�M.4�S5%CLv����L�;S�ڠ�� ɀ*^ДT���*��%��ue*��焘��v_#(壇v&�x}9�50�p/.�d����(�p#ȀH$"�-]��a�<�l&DlH���ݐ�I2����(�����|Y�KF�` ���J��ߟz�Kd�g3����ȸ�j��	��EF����g������6If�Q��RXGm1�B\�������(��L�7�l%�v �1��/Q���.E�3�W���V�����Î���E��i�P�4U
Шyd1�&���{�n����W+ń���ț�O�y�,�I���c�� 1��z��[G�?=�ˆ@��}qC��tQ7[�T��5F��(��jC�TwU,�m�=��j��0�"M�����d�&�lJ���-s�e*��A���կ~g���;��P.vѹ�k�K��d�C��o铧!Gw�n�ۙ���khK�L�v'wf������W38p�H�I�a��hIjY?i�-�}�b��?��r�ɩ9��#w��g��wF�`�Rudz$�Ew������;Eα�۷��5�b���d��y�kg�ᅺ��	�j��\�=�Д�N�r���ce��[��s�D᩿���p��v���������PWcҗ~O`�ԝ�� �a�d�>���&���4�m��f(8�(Ψ�6�U���2�t�e�C�Yk{1 SY�:���m#\B�Z����y���@ͦ�e������?2u���GrXF'�,�|:�u[�.6�:�V�U�~K��SO��5[Z��|^���V