��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$����r�/�/�Մ�����M�.,�W��˞��*t#�Ğ���W��OP�F���*k�=��l���˚N���g����r�]�K��4� hYc\���0�O�S@-� �S#
�h}R}��5sO �$��)�u�m-��P~e�R+]ă��&�}]�"�}�_-i�[�8V�?6x�:0�%n��k K��;��R�̌�J�4��f+S��A`=��Tcz��q�49���65`�zT{�f�B7h��z�n��76��>��$2���_Tp�'�ק�[DY�.kLvnP}S���+ʶ��F5�@�~�m���9�j���kJ���4������tMS��X��Ò�-�����z7qV���'�}�ā1hp*��n=��~���Mt�7$�>S�g�@�S��a�ڝ�.�,4,���`/�V�P]��	f��Z�jw��
�(�U����=�[~3D!�;�g��M��[�8�:W��t�Q��HZ�7嘊��ڵ�"?)�l� ��*���P4���+'j_��7叫��h�	�Z�ni���K�o|�c;�f��y+O:Z$�$p�[�y��B��6�i�úV��.�M�C\���&�L�r�u3kMVV4#����#�hMrX��2�z�#+-�Ykה~󲲦��PA<p���`&���YI?DM��^���N?LЃh�Z�!�`���O����ov�E$�=�!��a�rs1-�Mf��e����������|q7���r+8d�H,:��|zT�l,�y�`���D�[u�|M����O�PۦM£9 R�,�"?���C�H�"�B��k��R�,�S2�{�cu]������$�OX�wf�z�����J��P_����gq��e�^A����0z��B��O�F���x�Tg�*^ؤ]M�~�.���1E�Q�Y�e���[#�y�E��KŊL{�Ɛ���`��i!Zfs ���d�v����0�i�=\��A��?��� (��1_B�f�	�Ѻ+|n��y��Q4�]�aY�����*2�y%����>��������K������ �
�D��z�z��C�y�B����
_�U��hkF<�~x�ܕ�c�5�W���+u�k`�P�%b�L�nk��ӟ;v�a3bO��e�4Ҝ�FĒ�:�?\\t�Vޒ����Ƙ��|+�v�ϕ��َ� �]��IAx	6}��vF�k��ϋAi��9-`��P��3�����5:v�CG��#gb�)���k4�VW?��J�C��J\��k�ͅx=���#��:�o�R�e[h���bY���ޔ	ic0�0=��~b/B�]��x�Hu7ɖn��hﭥ/)��u��x����F��ۧ�XRr�:+��XT��";�Ci􈩳��]�x�3����8�Re����=a�+�aGIc:M2�WV*�K F�/�v�A��x�u��D�c�O�n��c��n��f��NdY=��8��
�\RΉ�����O�t���
���;�4F�M�1e�&�E��3�|:�^B�l�n7��T��M�j�����A��w#���*�Ő������/<!Cytv��ňl4�Aq�a�Ih�Ѱ��XS��#����m��G}��;��㋉�4��E��b��ߞ���p�m�yh7��[V�� .��t�*A4�}��G�̸L�վ~l��|Lז��_���S�ek��������=q0��_#�KaOL�����oY^�^-N���k	m(�{`V�NaJ՗(�n
��=���k�s:�-���171=/B%Ӱ�g���	���������<@����5�v��2�=-��!��Ϻ�$aYpB�!�e���22[���OR��Q���p�X��l�7�� �A�2�W�\�*U�'1Q22�%Dڤj�*��Tf�gDġ����o�0����O{W9���h����ö��t��6���0P0m��gAz'��@�78�;D�����+��nJL�sC۴~m��!�Z�a��}r�H�>)����.���G��|ѫ�����RtU9�mn�y�%�1I�5(˧}�NRx��xv�ۀ�s@������Y37 �m��8h�҄�J�F���%�+�����هȩF��.g�	���Y����3��N���啅�2;=�0��I�>�˃��Ҁ!���Φ ܔ�팻�O��Uh���2Sq��Sw<j~�Xp����z٭Z�z� v�;� ������0A��rH�����\1kꗍ��x�\��]f"�����LJ�y�K���_p���%:�}���Ư-�0@������p��obc8�_�Г�� ��5W�.��7�h����nd�,��H�ql��X��9���T y��^w;"�ܨk����J��.K^_��6'��G�p�,������4��~P=��)�
��=%7ls[�O~%K��f��'dH���{��փh�H�k5��
�C�����#�*"gJ	
��c�l� *}�@�M0$&^q�N|���k��O ��ʔi�Ɂg�&ı�f�.ɵ��n�5���'����U�A/ʦk�~��t4�Z���A����<'qWr܈c�aB���W����
t��KV�{q��� �;+��� �z'g���aeR�3f�;���ȏ�ऱJpk(>�BlY�o�W���iU]�j��E�����m	�}80��s_@��
�_� ��>���e��h��T@�F�$�Ҟ�iA�s[Ƭ�»�
R �������d�����K�1RrH�{�P��{J!���ko�"m#� kxr���h�ئGY�	��pe�a����=C�`�GԘ�z�����|�ݠ���QSB�}���{��o!h���g�iUR������$�}�C���I�[@����N���rn�d9}�ڷ�n��u{�,<~��|d�c����:p	���H��T��U>�Z��7�k�|�ɢ2N��Ȉ*�� �.g!�ݏ���(�d���q\���7�6]�5�3�%��轻ؑJ��8���>aNfY��ԇ��P�v�L�s����g)��wr&]�d�y2
����V��Fj0Y�ĳH�OMc}Yç.�;� ׀��(q8/h�C���?4�%8`2fs
�yM�˼XM�]ș� �r����8a�T�6��%j�Pt)���	K=ڰ�y}��?�
?�8��A_Y�P���J��O)q�c��D�H#ꁙ���v�B�PI�Fn�h�
�������/�Wy�,�{uC�l]ě ��B�}aʪ�usEB6�x�}Q�5��[̈7U���*��7���(4c1k��.�֕K�CR�qC
e3g�O���G��:W��w�y���75�}��`+�,?�A��K+�)8�K�xS�qyi��h�����I�P��)#v���u�<��">܌e�h?����.���/�q����Rw�i=�CA|g�U?��xk0��!`gh���9Q.;�'�es���m�b�zY���6d��ƛ����3����wx��]�@�6�8H�]���~�RZ�$�h��\-�~=�"q�U]ܽ�ȕm�'u]��Θ�[�ņ��>:|��QR��3���>~@èsr�T���?��� ��w�ڟ��m�0�P���Y�4�Y>kw��]Ń�^˥�k-J8x8�3�5cW;��K�Ո��-�4d�KQ� t%�Z:,�������$�u�p�˦��Ыf�L���g/h��6�B����uض����Yn��Ir���=�G�F��A��V=G8đ��rW�7�IB�Ox���t���@�� Tvyg�y��	��L%�s��_3��IzL:5�H�������7���������k��\ޒ�G�����۾Š�'�����z�j�K�1wA'���U���6�OC��&+ŁO�n���q7'��X���R��*�ߝ�"��;ȣ��<|JKv�Z���y��IOH�Aj�?xHy�r�=1���:�l��w�E�p��U2h�bu�
�f��\��|�T�,W~$Y��C�R�X�X�+&�ֹ�>)B���
t1Z�G#ɝ} ����g1��|�yّ����>ޖ#Q˘	�`>�R�T~5�(�z�a�C4Ql�u���o<�gY��L��J�Ǡ "����s���Μ��XBF�>�Ė*�K� �<-��]�E�(&ك1���M*@��>�'j?%��Js���g}��E�����XHFŕ�����}c�m�D(�L�^�aLф�Kc^�S�\�%��~	��s�	 )׃�� �>K���<���ٗ���/�/��;�i���`>�R@� ��+ä�Rr
�\������za� @��œ6"U�,pR0�/��ظ��Fƛ�Pc���d��V�ӣJa��{��p��<����Vة��r�`���=2��i64!R��H-�S,�cXp_����N���U�Vx��)!\v��!����*�z;��6�1����1!�?�~ޥ���~����t%���i_<�M�r�5A��TF~VFϼ�X��Y�X�=t����𨢸�� �_�>xD�����(Zί���Ng�Dv���`Åa�x�j���)����5l�G?m-9i���#�6Se?B�@ ���y_4�A�:����Q�~��9��(��z�� �l�F}CRDny�Qq4O�q��r�qUD�0.*ʷq�]Pe�� !#�[���h7��7����3E����b�Fֿ+.��$"KI�emй�idЀR�N[b���v�t i`������t��
�մo{E��>�T^#Vc��ԊW�8w��	?G�7K�h��iM;�t뛴&�ePd��2����a.q��52�� ��u"w�_��:�S�����	A�V�`Ӌ}�ig�`����&�G�Gr��5���Pj
�v7�n{q�|!�ܳ�v�y��������#�V3g?=Ctw�K��엷�K����?�ݾ���`(�u�b��/J�s^����k!VckI�Z��
�*qh�{A>z��}5)(��-#�����
�u�,���z�L�fsI<�LF������Ǽ+n����S6��P��~u���I(8Y�)���a(%q�DZsibY��5_�r��0�ƻ���ӗ'9L\�B���
��.LJ�G�^u!a&'��#Ob���9%�a�&�@�ʒ��\ڃ}#����B.����&��������Z;��--�`��~3j�a�Ͽ��:�J	�bb0k0�0y���Oҫ�����aM[��C���ﱐ�b��2Gm�P뽿���U�m��N��(����5� �����%?�d��>�B!��,l���iz��k��xD/�CX��N�3���wY��(�#�@I	]8s�"�%{I3��1z���HzI����9�w��'�>b�r��5¾���Qw��Ҿc>�v���S�8׌B�A*<a����4^�s@8������{���@��w��F�/���O�l���h86�Q�xַQ������@\���C�;�������T�B|x�$��O䱑��<%�(�3Eb��-��߮Kθul=�;�w�)�6
\�!+�H��,�_�S�î�S�⫤#���(�]ә�AI����z�N���A����Xj[�,^̐�PU�>z������Dp�����d�����!�ac0V9	/o�a.���;��!`919���V�	~�83�i�a#���������k�S:z�;�ɛ.OU�_ѺVF&�E��-�C����'�%�6���TxYd=*�+�4!�9!dC$pZт1j9���=hM�C�r�p��tf��ד����
���h,b�x�|vk�/��i:�º���M۟Y�r;�:��t��=) ���"jby�QߌvsΕV�'�U���M�I:�����d�o\�[��_�<Py\>�])j��+�1�G�B������G�?2�[�&���H O�Z��n�@�q��V�����%�W�~"_����L#t��VѸ�
(�k������|�9�q�Y�K;���}c����P�����6ir�P�h/?��;��x���^�ښ4��mƕꡮ��p+q�m{)��G���7+:`�+V�g>G�e�ՖɦѶ_�hN��S�%/zΉ�4�ÃS K��|d�:�kpˈGos�OG�0>{���8�d{��G�!7�||<�tM�Y�SE5N��OYy��@�3���j�`@���^�3 �4�Z��9��f}�B?��Z�~��}�w:_�#
���t�#��8ľk��3����N��;����x8.H�2$�=��!8&�f�����$>g����K����xU�$k��0��I-�:���ϘrV*�R�}��+�ڑ>�u3T0A�߄bN�=m��k�$��Bn��h#G�@�/��r�m�1QT��:�_���z���W��\Om8�b����ԏɦ��*H����q ����n=���\�JH��bW]q�S����3|��ԛ⛔�\�A��W�,'��1�.�P!ZC2!�&�|�h��-��q����u�}.�� _�l �h�3,(&,�Y�թ��/e�8��:�qd'�?`ܕ �^�%��^?���4�<��8�_��D����(���I�&c��	��M��e��PG&�\Q�N� V[a�� ��T��K�f��l���p[u��9��0T@�B��lg���e�b7�m�,�T������HM�Y��ۋz��^h�_Fok���;6�.�L{ĝ?�c��E�GIV�%����,���["�v��vj�K����R$]��7�b����|��#��jH7�'�Y�:���8¤�(�"<��ج�����	�vs]�-P�$��\���?!Bw��,���v&z�;��?!��h�A��:s�MB�|��W�*s	�6H�¸ ��a��B+��g�;��ޯ�.��Hp`4ȅi���l���xG<}�*�7.�L~�^�xO��+O��y�\_z�����M�W��p΂K���r.f]M��xW��FG�;�c�I���f}#��w����Pe�z��q���5I�L���L�U�h�H��ʜc��~�.D�q����4�@���+��h��3S��gR�֗$���X+�gve+S�lC0]k_[_���(��5�E�[����.��{��YZ'5��9_C�ٗ�}���u���]�Q]㡎�jC���>�Ծ��A͠�S���7����-�%�]lp`�i�=.|Z�S+�8H�-�&��14�}�R�M��ڐ�"%�h��]*��|�w#�������J�gL�ӯ�HR���ˋ5b���4�D@���)�85�_�P~�q[�uE˯��j������r@�7�s�>����~����f3��1<��2�j���]}QZRJZ�W�\�2&�{�:t/���w?,�&B�4i桄�l��B��ctF�O�-�g C��;'�trһB$QGҖdS�ҏ�+Ӊ�4�b5����~p��a���әt !�}�^���X\�v�3�G:;:6cG�����/�/a뻽Q>�2���.4v�;B���GUc-�	7H�
�d�qC�'${ C�Ɗ��(�P�VmMg�t�Ϟ�`E�[cO �i�$�QF�nEK�{֜n��{u��/j2���U.��N��t��)Yk:�)��VV��i)���O������a-�B��^�}�ߤ�	��5��ksz��t�t��uV���(��}����^��̏}�Ql��M�-�sV���	���y��6���W>��w��X:��� "R*��!Q��n>tV;�/��2���h����hz��?�;^��n�:p��͔��{R�GA�}C�	vi}���mX���%�_�>@���(�۫��7�S�2��Ik����0D��( ���;�����SP�o ���Ӫ%�ٲ �ĸ\͙�j���ی��W!� r��o�&��`���Z6�5ˀ�t<�2V�;*�����0�	ON�5H���_�j!����M�:u�RΆ <�?�^�k����蛦 TA��L4�$�i�{�&%��߈	�������=˳���r3���H��I�D!#{�T�@@���"�zb`o�����`����nԩ{��ԇЉ��>[L���� ��/�˽ނL��r'Q������=�K_��/3c����?H65�,_���������KOA&/@�V2Y��Z~�J��EV=ۖѵ$��逝�{�:?YM-J����#P�*�'�Cq�ޣ�1�-�AF�1�\+�:3�am0_?���5���	f����q��?������x��}5|��5��zuL�ly
�'�3��E��&�I�8��rk�����ʝ�yv�/��)}�F�{�[ OW��%����
nN����>v�5o�ԽE�h�Hk�6��l0�)����N0�jv438)�r�)rb x�-gD�����P䀳�1��V۱�`/��s�
�(%���t�є2/���uWoy%�T��?9m��a�.�Tf�
��Ӕ����i����ԡ<
t-
"�S�O>��"�`�0���9CPu>�e�&��â��
��U_�u��t���G��W`2������$X�S�ļ?�2F'�����*�����&@��zm*"��4nXy��z���`�����K$��ʅ��� ��[v^y���u0�*
�Mw�7+çӌ����uw]K'�|�n�G��e�ԡ%�%��8�.�et�t#� J�t�C�;1	1���ZӮ��>	�M�hyf��G#H�q�ZϣrSO|ɳ_]�h��3�`��<�NxAZ��L6x��@Þc{�(*s�L���JR�]��V�i�Eq�Y��Y�hC~n�f�(eo�n	؅��Y��!�u��b�J26��!ݼ�=] M�%�����[�ۏ�>��Vy0+�Ki&�>٦@kAS	�}�4�rW='x�lL^_*���J�.���x��)=�ZpuM��=`�C\�9RO�R��V�\^�U���п+�i߃��N�iUr��
m)	��l��� "��(��c�_`u����Vr�E�ޒLT�U�&�R�\ǔf�Բ~A�I94VGm��R�fpeb��a���ꃧ��m�
gB�M���:k38����Ǐ��I6n�PN��Q*>y@3�B��\��Kbҷ%�)�D���x�$E��_9qB|�`}Xx�+�c$�Y]z����{Pz�{��t�~� �뚁���X��z\B��]�]2gۇB�1'a�Wg���)�D�� H�j�NÑO���Yϙ��F3zx���ۑ�/W�V#?�`{�Y�i��
YKzм��S��C�!/F�M:�OvE����d-�1��H�����ـT� R�Y�dJ��
$XA �^l��OHE�E�ɺB��]2�����SvռX��#�n�$:t�-k��As#O��эGf�m3gi��Ji	��"�E��ιRf0G-��E<9h0��4��#���-��W
�J�k�?hu�@�)�?�@z�!	o�;/���	��aN��u9�|ÆU���X޴"Szm*�;tM5����5�Mk�7,�:b���j�����&�2J�I9,�~��W����HvN����ء9��u�ƹ��&�kIД)�n�x�"0 �@��S��m����p��CKz�ZQ�������Y��ŧ	�"gU�y@��̬���=A�¾�1�F�l6����m�D�^�o��S��^�Q��d��Wk�x��>��m]����ġ~T�� ��vu|w˝�l�G�&.�Gzr(C$bފF̶��^p���-a^5�J���Y�=��]�b=ֺ8u�E�#��/��Vi 5fne�6����9�Z�]83�f��^��-���j�6�zOG^И��e�w�k��\�̑_U�q�r�����8#/�`�o��f\��p!Wbm~�m�q�'�=R+[e0�'����&^��U��A߶����"�����譍�/"�k��}m��.Nb��&T�����f1����vX�f_��RO�$��������q9����e,�͊B�Z���HY$
w�
�H��O�N�&ġ�2Pl���p����!�d�/!�T�!�u��9��������Kp#�+��u��Jve�C����� D��}�Iv��$��\��f%��t,�7ol�&���
�����f90&��lܞ���ɥ��'����
���v���V��Mr��n�T4f �K�uCV�P�s���P	��,ݲ�]KI��Z��
� �밑���.��[�<���`|4ú�b�tO�����-���"��d����	��F}ͮ[x�V8�DC�-�i� Q����[�ҟ��A���U��ag�ڜ$b�Q^X���%f��n����&]4~�&ξݝ���f��ʦ���A�*�В�Le�din�	J�2ץBW
40a�oK0�ƨ*�q�l�6�f±L)�]V�(�����ĿeΦ mW#rT��	4.>�Ww+.��tR�-�!�#S�[=P�}�J�~�뫓�]%8��I�(Qm��"m�����Ib��7�a���m{XlB�5��!���d >��?�IaI�^;�F�mM�'���z"5��n�g�Ue�xK�z���$IH&�p���I�Ǧxl�����k��<�~�;���k7g��YU��V�F!�+�/2^FNܡ��=B�`G7%��m\�&����߂W����d?��mm��D$3$xVg%v,r��@�C�K�f��/V��I��� v}�
B�w�Qz���63C1nD�3]��SF3}�_�(xXW��=I�Y�e8Z�5�f�U\����D��v�M3�&�_�\X�ܽ�]08Fz����q���_alKɬ�@�l����~t��X�T�����S��{�G
f���Z�d:�7����>������C���/�Q|\��H��m!_p����9�
�%��|�.5��LU1w%���Y��@Ԟ�>ܙ""X�;��3?��Jݰ�p�b�@^᳘M`���C�r�y�Y����Tm��6�[
$\*h�D�3;-QM��2���'7��ۘ���H�a�(ǿa5�;��B��$2UN=�T7�j� -R���j&l�z9J��E&@.�c����s��˥��~���}����nF(�@��@���|�Ɣ�O~�����Y�3�&"�W3P2���ui�l��&׷0�c�s��x#)��9�O�I>ϟG�n���"E���b\Rf� �%�p�ڙ��ǫk^;s~�x���Yv���i5��L�L �B���R�#u| U�:����un�z��/��w}D���j���z�K��N�	��;�����)4&���=wϹD�����2ؕ���6�+����$=~ۮ���ʁ.q:�cC��}���sw�Fh.��!��K�L�vT��[��ii��&�㬙�
n�O��	?���Z�
��4��^�+��}���muo�2��`v�b�q3Ч,�S�}C��M�`�Q�m:y�X=�����)Iz.���L����{am�c&f�?�ֳ6�9+=_�)W}�]Q�S�����aW� E���GF�*�����O��˸��{"�G�9�C=A�Xe��@��ö��mXMb7Ŝ�1�0M�ZA��f�ǫ�/n]���5V��~�5�F��^5�g3%�5ڑ�RŹ ������\=�č�"Uk%2�"�{�)S���"-b�WDNjr�����J���+ ��'�?Y)�E�C�v� W?�i�O�6�k #�b6�WZ K$����<�;�t���?3P~+Le/�K|��z{0 Âe<po��鸳g�|
�}��y��W�3��x@�Ʈ�D3��yWu�u�8���⦂)��jc^L++��e1Y���/���"v{):ė�;'�)�oZ����$���K�i���j�C�J�3Ϲ�4� �sr
<=M�@���<�X�`[Ї�+C<:T�Bx<"k�z����+]�-�O��j��g;9O����w�8�p���֖2�p�p�yC!�x���ty ��;�
�>'<z��C'���r����Y���2�z������